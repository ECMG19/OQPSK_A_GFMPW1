magic
tech gf180mcuD
magscale 1 5
timestamp 1701968756
<< obsm1 >>
rect 672 1538 29288 28321
<< metal2 >>
rect 2688 29600 2744 30000
rect 3024 29600 3080 30000
rect 3696 29600 3752 30000
rect 4368 29600 4424 30000
rect 4704 29600 4760 30000
rect 5376 29600 5432 30000
rect 5712 29600 5768 30000
rect 15456 29600 15512 30000
rect 20496 29600 20552 30000
rect 22848 29600 22904 30000
rect 26208 29600 26264 30000
rect 27216 29600 27272 30000
rect 27552 29600 27608 30000
rect 2352 0 2408 400
rect 4704 0 4760 400
rect 14448 0 14504 400
rect 21168 0 21224 400
rect 21840 0 21896 400
rect 23184 0 23240 400
rect 25200 0 25256 400
rect 25536 0 25592 400
rect 26208 0 26264 400
<< obsm2 >>
rect 854 29570 2658 29600
rect 2774 29570 2994 29600
rect 3110 29570 3666 29600
rect 3782 29570 4338 29600
rect 4454 29570 4674 29600
rect 4790 29570 5346 29600
rect 5462 29570 5682 29600
rect 5798 29570 15426 29600
rect 15542 29570 20466 29600
rect 20582 29570 22818 29600
rect 22934 29570 26178 29600
rect 26294 29570 27186 29600
rect 27302 29570 27522 29600
rect 27638 29570 29162 29600
rect 854 430 29162 29570
rect 854 400 2322 430
rect 2438 400 4674 430
rect 4790 400 14418 430
rect 14534 400 21138 430
rect 21254 400 21810 430
rect 21926 400 23154 430
rect 23270 400 25170 430
rect 25286 400 25506 430
rect 25622 400 26178 430
rect 26294 400 29162 430
<< metal3 >>
rect 0 27216 400 27272
rect 29600 26544 30000 26600
rect 0 25536 400 25592
rect 29600 25200 30000 25256
rect 29600 24864 30000 24920
rect 0 24192 400 24248
rect 0 23856 400 23912
rect 29600 23520 30000 23576
rect 29600 22176 30000 22232
rect 29600 21504 30000 21560
rect 0 21168 400 21224
rect 0 20496 400 20552
rect 29600 20160 30000 20216
rect 0 19488 400 19544
rect 29600 18816 30000 18872
rect 0 18480 400 18536
rect 0 18144 400 18200
rect 0 17808 400 17864
rect 29600 17808 30000 17864
rect 0 17472 400 17528
rect 29600 17472 30000 17528
rect 0 16800 400 16856
rect 0 16464 400 16520
rect 29600 16464 30000 16520
rect 0 15792 400 15848
rect 0 15456 400 15512
rect 0 15120 400 15176
rect 29600 15120 30000 15176
rect 0 14784 400 14840
rect 0 14448 400 14504
rect 0 14112 400 14168
rect 29600 14112 30000 14168
rect 0 13776 400 13832
rect 0 13440 400 13496
rect 29600 13104 30000 13160
rect 0 12768 400 12824
rect 29600 12768 30000 12824
rect 29600 12432 30000 12488
rect 0 12096 400 12152
rect 29600 11760 30000 11816
rect 29600 11088 30000 11144
rect 29600 10752 30000 10808
rect 0 10416 400 10472
rect 29600 9744 30000 9800
rect 29600 9408 30000 9464
rect 29600 9072 30000 9128
rect 0 8736 400 8792
rect 29600 8400 30000 8456
rect 29600 8064 30000 8120
rect 29600 7728 30000 7784
rect 29600 6720 30000 6776
rect 29600 6048 30000 6104
rect 29600 5712 30000 5768
rect 29600 5376 30000 5432
rect 29600 5040 30000 5096
rect 29600 4704 30000 4760
rect 29600 4368 30000 4424
rect 29600 4032 30000 4088
<< obsm3 >>
rect 400 27302 29666 28938
rect 430 27186 29666 27302
rect 400 26630 29666 27186
rect 400 26514 29570 26630
rect 400 25622 29666 26514
rect 430 25506 29666 25622
rect 400 25286 29666 25506
rect 400 25170 29570 25286
rect 400 24950 29666 25170
rect 400 24834 29570 24950
rect 400 24278 29666 24834
rect 430 24162 29666 24278
rect 400 23942 29666 24162
rect 430 23826 29666 23942
rect 400 23606 29666 23826
rect 400 23490 29570 23606
rect 400 22262 29666 23490
rect 400 22146 29570 22262
rect 400 21590 29666 22146
rect 400 21474 29570 21590
rect 400 21254 29666 21474
rect 430 21138 29666 21254
rect 400 20582 29666 21138
rect 430 20466 29666 20582
rect 400 20246 29666 20466
rect 400 20130 29570 20246
rect 400 19574 29666 20130
rect 430 19458 29666 19574
rect 400 18902 29666 19458
rect 400 18786 29570 18902
rect 400 18566 29666 18786
rect 430 18450 29666 18566
rect 400 18230 29666 18450
rect 430 18114 29666 18230
rect 400 17894 29666 18114
rect 430 17778 29570 17894
rect 400 17558 29666 17778
rect 430 17442 29570 17558
rect 400 16886 29666 17442
rect 430 16770 29666 16886
rect 400 16550 29666 16770
rect 430 16434 29570 16550
rect 400 15878 29666 16434
rect 430 15762 29666 15878
rect 400 15542 29666 15762
rect 430 15426 29666 15542
rect 400 15206 29666 15426
rect 430 15090 29570 15206
rect 400 14870 29666 15090
rect 430 14754 29666 14870
rect 400 14534 29666 14754
rect 430 14418 29666 14534
rect 400 14198 29666 14418
rect 430 14082 29570 14198
rect 400 13862 29666 14082
rect 430 13746 29666 13862
rect 400 13526 29666 13746
rect 430 13410 29666 13526
rect 400 13190 29666 13410
rect 400 13074 29570 13190
rect 400 12854 29666 13074
rect 430 12738 29570 12854
rect 400 12518 29666 12738
rect 400 12402 29570 12518
rect 400 12182 29666 12402
rect 430 12066 29666 12182
rect 400 11846 29666 12066
rect 400 11730 29570 11846
rect 400 11174 29666 11730
rect 400 11058 29570 11174
rect 400 10838 29666 11058
rect 400 10722 29570 10838
rect 400 10502 29666 10722
rect 430 10386 29666 10502
rect 400 9830 29666 10386
rect 400 9714 29570 9830
rect 400 9494 29666 9714
rect 400 9378 29570 9494
rect 400 9158 29666 9378
rect 400 9042 29570 9158
rect 400 8822 29666 9042
rect 430 8706 29666 8822
rect 400 8486 29666 8706
rect 400 8370 29570 8486
rect 400 8150 29666 8370
rect 400 8034 29570 8150
rect 400 7814 29666 8034
rect 400 7698 29570 7814
rect 400 6806 29666 7698
rect 400 6690 29570 6806
rect 400 6134 29666 6690
rect 400 6018 29570 6134
rect 400 5798 29666 6018
rect 400 5682 29570 5798
rect 400 5462 29666 5682
rect 400 5346 29570 5462
rect 400 5126 29666 5346
rect 400 5010 29570 5126
rect 400 4790 29666 5010
rect 400 4674 29570 4790
rect 400 4454 29666 4674
rect 400 4338 29570 4454
rect 400 4118 29666 4338
rect 400 4002 29570 4118
rect 400 686 29666 4002
<< metal4 >>
rect 2224 1538 2384 28254
rect 9904 1538 10064 28254
rect 17584 1538 17744 28254
rect 25264 1538 25424 28254
<< obsm4 >>
rect 3430 28284 23282 28943
rect 3430 1508 9874 28284
rect 10094 1508 17554 28284
rect 17774 1508 23282 28284
rect 3430 681 23282 1508
<< labels >>
rlabel metal3 s 29600 15120 30000 15176 6 BitIn
port 1 nsew signal input
rlabel metal3 s 0 16800 400 16856 6 CLK
port 2 nsew signal input
rlabel metal3 s 0 15456 400 15512 6 EN
port 3 nsew signal input
rlabel metal3 s 29600 12432 30000 12488 6 I[0]
port 4 nsew signal output
rlabel metal2 s 23184 0 23240 400 6 I[10]
port 5 nsew signal output
rlabel metal2 s 21840 0 21896 400 6 I[11]
port 6 nsew signal output
rlabel metal2 s 21168 0 21224 400 6 I[12]
port 7 nsew signal output
rlabel metal3 s 29600 11760 30000 11816 6 I[1]
port 8 nsew signal output
rlabel metal3 s 29600 10752 30000 10808 6 I[2]
port 9 nsew signal output
rlabel metal3 s 29600 9072 30000 9128 6 I[3]
port 10 nsew signal output
rlabel metal3 s 29600 8400 30000 8456 6 I[4]
port 11 nsew signal output
rlabel metal3 s 29600 7728 30000 7784 6 I[5]
port 12 nsew signal output
rlabel metal3 s 29600 5712 30000 5768 6 I[6]
port 13 nsew signal output
rlabel metal3 s 29600 4368 30000 4424 6 I[7]
port 14 nsew signal output
rlabel metal2 s 25536 0 25592 400 6 I[8]
port 15 nsew signal output
rlabel metal2 s 25200 0 25256 400 6 I[9]
port 16 nsew signal output
rlabel metal2 s 20496 29600 20552 30000 6 Q[0]
port 17 nsew signal output
rlabel metal3 s 29600 17472 30000 17528 6 Q[10]
port 18 nsew signal output
rlabel metal3 s 29600 16464 30000 16520 6 Q[11]
port 19 nsew signal output
rlabel metal3 s 29600 17808 30000 17864 6 Q[12]
port 20 nsew signal output
rlabel metal2 s 22848 29600 22904 30000 6 Q[1]
port 21 nsew signal output
rlabel metal2 s 26208 29600 26264 30000 6 Q[2]
port 22 nsew signal output
rlabel metal3 s 29600 26544 30000 26600 6 Q[3]
port 23 nsew signal output
rlabel metal3 s 29600 25200 30000 25256 6 Q[4]
port 24 nsew signal output
rlabel metal3 s 29600 24864 30000 24920 6 Q[5]
port 25 nsew signal output
rlabel metal3 s 29600 22176 30000 22232 6 Q[6]
port 26 nsew signal output
rlabel metal3 s 29600 21504 30000 21560 6 Q[7]
port 27 nsew signal output
rlabel metal3 s 29600 20160 30000 20216 6 Q[8]
port 28 nsew signal output
rlabel metal3 s 29600 18816 30000 18872 6 Q[9]
port 29 nsew signal output
rlabel metal3 s 0 16464 400 16520 6 RST
port 30 nsew signal input
rlabel metal3 s 0 13776 400 13832 6 addI[0]
port 31 nsew signal output
rlabel metal3 s 0 14112 400 14168 6 addI[1]
port 32 nsew signal output
rlabel metal3 s 0 14784 400 14840 6 addI[2]
port 33 nsew signal output
rlabel metal3 s 0 14448 400 14504 6 addI[3]
port 34 nsew signal output
rlabel metal3 s 0 15120 400 15176 6 addI[4]
port 35 nsew signal output
rlabel metal2 s 14448 0 14504 400 6 addI[5]
port 36 nsew signal output
rlabel metal3 s 0 17472 400 17528 6 addQ[0]
port 37 nsew signal output
rlabel metal3 s 0 18144 400 18200 6 addQ[1]
port 38 nsew signal output
rlabel metal3 s 0 23856 400 23912 6 addQ[2]
port 39 nsew signal output
rlabel metal3 s 0 24192 400 24248 6 addQ[3]
port 40 nsew signal output
rlabel metal3 s 0 27216 400 27272 6 addQ[4]
port 41 nsew signal output
rlabel metal2 s 15456 29600 15512 30000 6 addQ[5]
port 42 nsew signal output
rlabel metal3 s 0 12096 400 12152 6 io_oeb[0]
port 43 nsew signal output
rlabel metal3 s 29600 14112 30000 14168 6 io_oeb[10]
port 44 nsew signal output
rlabel metal3 s 29600 5040 30000 5096 6 io_oeb[11]
port 45 nsew signal output
rlabel metal2 s 3024 29600 3080 30000 6 io_oeb[12]
port 46 nsew signal output
rlabel metal3 s 0 19488 400 19544 6 io_oeb[13]
port 47 nsew signal output
rlabel metal3 s 29600 9408 30000 9464 6 io_oeb[14]
port 48 nsew signal output
rlabel metal3 s 0 8736 400 8792 6 io_oeb[15]
port 49 nsew signal output
rlabel metal2 s 5376 29600 5432 30000 6 io_oeb[16]
port 50 nsew signal output
rlabel metal3 s 0 25536 400 25592 6 io_oeb[17]
port 51 nsew signal output
rlabel metal3 s 29600 13104 30000 13160 6 io_oeb[18]
port 52 nsew signal output
rlabel metal3 s 29600 12768 30000 12824 6 io_oeb[19]
port 53 nsew signal output
rlabel metal3 s 0 20496 400 20552 6 io_oeb[1]
port 54 nsew signal output
rlabel metal3 s 0 17808 400 17864 6 io_oeb[20]
port 55 nsew signal output
rlabel metal3 s 0 15792 400 15848 6 io_oeb[21]
port 56 nsew signal output
rlabel metal3 s 29600 4704 30000 4760 6 io_oeb[22]
port 57 nsew signal output
rlabel metal3 s 29600 8064 30000 8120 6 io_oeb[23]
port 58 nsew signal output
rlabel metal3 s 29600 11088 30000 11144 6 io_oeb[24]
port 59 nsew signal output
rlabel metal2 s 27216 29600 27272 30000 6 io_oeb[25]
port 60 nsew signal output
rlabel metal2 s 4704 0 4760 400 6 io_oeb[26]
port 61 nsew signal output
rlabel metal3 s 0 10416 400 10472 6 io_oeb[27]
port 62 nsew signal output
rlabel metal2 s 4704 29600 4760 30000 6 io_oeb[28]
port 63 nsew signal output
rlabel metal3 s 29600 4032 30000 4088 6 io_oeb[29]
port 64 nsew signal output
rlabel metal3 s 0 12768 400 12824 6 io_oeb[2]
port 65 nsew signal output
rlabel metal2 s 26208 0 26264 400 6 io_oeb[30]
port 66 nsew signal output
rlabel metal3 s 29600 9744 30000 9800 6 io_oeb[31]
port 67 nsew signal output
rlabel metal2 s 27552 29600 27608 30000 6 io_oeb[32]
port 68 nsew signal output
rlabel metal2 s 2352 0 2408 400 6 io_oeb[33]
port 69 nsew signal output
rlabel metal3 s 0 13440 400 13496 6 io_oeb[34]
port 70 nsew signal output
rlabel metal3 s 29600 6048 30000 6104 6 io_oeb[35]
port 71 nsew signal output
rlabel metal2 s 5712 29600 5768 30000 6 io_oeb[36]
port 72 nsew signal output
rlabel metal2 s 2688 29600 2744 30000 6 io_oeb[37]
port 73 nsew signal output
rlabel metal3 s 0 21168 400 21224 6 io_oeb[3]
port 74 nsew signal output
rlabel metal3 s 29600 5376 30000 5432 6 io_oeb[4]
port 75 nsew signal output
rlabel metal2 s 4368 29600 4424 30000 6 io_oeb[5]
port 76 nsew signal output
rlabel metal3 s 0 18480 400 18536 6 io_oeb[6]
port 77 nsew signal output
rlabel metal3 s 29600 23520 30000 23576 6 io_oeb[7]
port 78 nsew signal output
rlabel metal3 s 29600 6720 30000 6776 6 io_oeb[8]
port 79 nsew signal output
rlabel metal2 s 3696 29600 3752 30000 6 io_oeb[9]
port 80 nsew signal output
rlabel metal4 s 2224 1538 2384 28254 6 vdd
port 81 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 28254 6 vdd
port 81 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 28254 6 vss
port 82 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 28254 6 vss
port 82 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 30000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3160628
string GDS_FILE /home/emmascorro/Escritorio/Proyectos_caravel/OQPSK_S_GFMPW1/openlane/OQPSK_S_GFMPW1/runs/23_12_07_11_03/results/signoff/OQPSK_PS_RCOSINE2.magic.gds
string GDS_START 481472
<< end >>

