magic
tech gf180mcuD
magscale 1 10
timestamp 1701968754
<< metal1 >>
rect 54450 56590 54462 56642
rect 54514 56639 54526 56642
rect 55010 56639 55022 56642
rect 54514 56593 55022 56639
rect 54514 56590 54526 56593
rect 55010 56590 55022 56593
rect 55074 56590 55086 56642
rect 1344 56474 58576 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 58576 56474
rect 1344 56388 58576 56422
rect 5630 56306 5682 56318
rect 5630 56242 5682 56254
rect 6302 56306 6354 56318
rect 6302 56242 6354 56254
rect 7646 56306 7698 56318
rect 7646 56242 7698 56254
rect 9662 56306 9714 56318
rect 9662 56242 9714 56254
rect 11006 56306 11058 56318
rect 11006 56242 11058 56254
rect 11678 56306 11730 56318
rect 11678 56242 11730 56254
rect 18286 56306 18338 56318
rect 18286 56242 18338 56254
rect 21086 56306 21138 56318
rect 27022 56306 27074 56318
rect 23314 56254 23326 56306
rect 23378 56254 23390 56306
rect 21086 56242 21138 56254
rect 27022 56242 27074 56254
rect 48414 56306 48466 56318
rect 48414 56242 48466 56254
rect 55022 56306 55074 56318
rect 55022 56242 55074 56254
rect 55470 56306 55522 56318
rect 55470 56242 55522 56254
rect 13806 56194 13858 56206
rect 13806 56130 13858 56142
rect 19182 56194 19234 56206
rect 19182 56130 19234 56142
rect 21870 56194 21922 56206
rect 25566 56194 25618 56206
rect 24658 56142 24670 56194
rect 24722 56142 24734 56194
rect 21870 56130 21922 56142
rect 25566 56130 25618 56142
rect 28478 56194 28530 56206
rect 28478 56130 28530 56142
rect 28702 56194 28754 56206
rect 28702 56130 28754 56142
rect 37438 56194 37490 56206
rect 37438 56130 37490 56142
rect 19070 56082 19122 56094
rect 30718 56082 30770 56094
rect 36990 56082 37042 56094
rect 19730 56030 19742 56082
rect 19794 56030 19806 56082
rect 21298 56030 21310 56082
rect 21362 56030 21374 56082
rect 24546 56030 24558 56082
rect 24610 56030 24622 56082
rect 31490 56030 31502 56082
rect 31554 56030 31566 56082
rect 34290 56030 34302 56082
rect 34354 56030 34366 56082
rect 42578 56030 42590 56082
rect 42642 56030 42654 56082
rect 47394 56030 47406 56082
rect 47458 56030 47470 56082
rect 54002 56030 54014 56082
rect 54066 56030 54078 56082
rect 19070 56018 19122 56030
rect 30718 56018 30770 56030
rect 36990 56018 37042 56030
rect 8766 55970 8818 55982
rect 8766 55906 8818 55918
rect 14142 55970 14194 55982
rect 14142 55906 14194 55918
rect 14702 55970 14754 55982
rect 14702 55906 14754 55918
rect 15150 55970 15202 55982
rect 15150 55906 15202 55918
rect 15598 55970 15650 55982
rect 15598 55906 15650 55918
rect 16046 55970 16098 55982
rect 16046 55906 16098 55918
rect 16494 55970 16546 55982
rect 16494 55906 16546 55918
rect 17502 55970 17554 55982
rect 17502 55906 17554 55918
rect 17950 55970 18002 55982
rect 17950 55906 18002 55918
rect 18846 55970 18898 55982
rect 23102 55970 23154 55982
rect 20066 55918 20078 55970
rect 20130 55918 20142 55970
rect 18846 55906 18898 55918
rect 23102 55906 23154 55918
rect 26126 55970 26178 55982
rect 26126 55906 26178 55918
rect 26798 55970 26850 55982
rect 26798 55906 26850 55918
rect 27582 55970 27634 55982
rect 27582 55906 27634 55918
rect 29598 55970 29650 55982
rect 29598 55906 29650 55918
rect 30158 55970 30210 55982
rect 30158 55906 30210 55918
rect 31054 55970 31106 55982
rect 31054 55906 31106 55918
rect 32398 55970 32450 55982
rect 32398 55906 32450 55918
rect 35310 55970 35362 55982
rect 35310 55906 35362 55918
rect 36094 55970 36146 55982
rect 36094 55906 36146 55918
rect 36542 55970 36594 55982
rect 41010 55918 41022 55970
rect 41074 55918 41086 55970
rect 52434 55918 52446 55970
rect 52498 55918 52510 55970
rect 36542 55906 36594 55918
rect 19182 55858 19234 55870
rect 15138 55806 15150 55858
rect 15202 55855 15214 55858
rect 16482 55855 16494 55858
rect 15202 55809 16494 55855
rect 15202 55806 15214 55809
rect 16482 55806 16494 55809
rect 16546 55806 16558 55858
rect 19182 55794 19234 55806
rect 24670 55858 24722 55870
rect 24670 55794 24722 55806
rect 28366 55858 28418 55870
rect 28366 55794 28418 55806
rect 1344 55690 58576 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 58576 55690
rect 1344 55604 58576 55638
rect 18062 55522 18114 55534
rect 18062 55458 18114 55470
rect 19070 55522 19122 55534
rect 19070 55458 19122 55470
rect 1934 55410 1986 55422
rect 1934 55346 1986 55358
rect 14142 55410 14194 55422
rect 14142 55346 14194 55358
rect 17838 55410 17890 55422
rect 24334 55410 24386 55422
rect 19618 55358 19630 55410
rect 19682 55358 19694 55410
rect 22642 55358 22654 55410
rect 22706 55358 22718 55410
rect 26786 55358 26798 55410
rect 26850 55358 26862 55410
rect 30258 55358 30270 55410
rect 30322 55358 30334 55410
rect 37874 55358 37886 55410
rect 37938 55358 37950 55410
rect 47954 55358 47966 55410
rect 48018 55358 48030 55410
rect 17838 55346 17890 55358
rect 24334 55346 24386 55358
rect 15934 55298 15986 55310
rect 4162 55246 4174 55298
rect 4226 55246 4238 55298
rect 15934 55234 15986 55246
rect 18734 55298 18786 55310
rect 23998 55298 24050 55310
rect 28254 55298 28306 55310
rect 31166 55298 31218 55310
rect 19058 55246 19070 55298
rect 19122 55246 19134 55298
rect 20738 55246 20750 55298
rect 20802 55246 20814 55298
rect 21746 55246 21758 55298
rect 21810 55246 21822 55298
rect 23762 55246 23774 55298
rect 23826 55246 23838 55298
rect 26674 55246 26686 55298
rect 26738 55246 26750 55298
rect 29810 55246 29822 55298
rect 29874 55246 29886 55298
rect 18734 55234 18786 55246
rect 23998 55234 24050 55246
rect 28254 55234 28306 55246
rect 31166 55234 31218 55246
rect 32174 55298 32226 55310
rect 32174 55234 32226 55246
rect 33854 55298 33906 55310
rect 33854 55234 33906 55246
rect 34414 55298 34466 55310
rect 36206 55298 36258 55310
rect 40910 55298 40962 55310
rect 44046 55298 44098 55310
rect 35970 55246 35982 55298
rect 36034 55246 36046 55298
rect 37538 55246 37550 55298
rect 37602 55246 37614 55298
rect 40338 55246 40350 55298
rect 40402 55246 40414 55298
rect 43362 55246 43374 55298
rect 43426 55246 43438 55298
rect 43810 55246 43822 55298
rect 43874 55246 43886 55298
rect 34414 55234 34466 55246
rect 36206 55234 36258 55246
rect 40910 55234 40962 55246
rect 44046 55234 44098 55246
rect 44942 55298 44994 55310
rect 51214 55298 51266 55310
rect 45266 55246 45278 55298
rect 45330 55246 45342 55298
rect 51426 55246 51438 55298
rect 51490 55246 51502 55298
rect 44942 55234 44994 55246
rect 51214 55234 51266 55246
rect 15038 55186 15090 55198
rect 15038 55122 15090 55134
rect 15374 55186 15426 55198
rect 15374 55122 15426 55134
rect 16494 55186 16546 55198
rect 16494 55122 16546 55134
rect 17390 55186 17442 55198
rect 17390 55122 17442 55134
rect 22206 55186 22258 55198
rect 22206 55122 22258 55134
rect 27918 55186 27970 55198
rect 27918 55122 27970 55134
rect 28478 55186 28530 55198
rect 28478 55122 28530 55134
rect 32734 55186 32786 55198
rect 32734 55122 32786 55134
rect 33070 55186 33122 55198
rect 33070 55122 33122 55134
rect 34862 55186 34914 55198
rect 34862 55122 34914 55134
rect 36430 55186 36482 55198
rect 36430 55122 36482 55134
rect 37214 55186 37266 55198
rect 37214 55122 37266 55134
rect 38222 55186 38274 55198
rect 38222 55122 38274 55134
rect 41022 55186 41074 55198
rect 41022 55122 41074 55134
rect 41358 55186 41410 55198
rect 41358 55122 41410 55134
rect 41694 55186 41746 55198
rect 41694 55122 41746 55134
rect 42478 55186 42530 55198
rect 42478 55122 42530 55134
rect 42702 55186 42754 55198
rect 42702 55122 42754 55134
rect 45838 55186 45890 55198
rect 45838 55122 45890 55134
rect 46174 55186 46226 55198
rect 46174 55122 46226 55134
rect 46510 55186 46562 55198
rect 49870 55186 49922 55198
rect 48178 55134 48190 55186
rect 48242 55134 48254 55186
rect 46510 55122 46562 55134
rect 49870 55122 49922 55134
rect 52110 55186 52162 55198
rect 52110 55122 52162 55134
rect 52670 55186 52722 55198
rect 52670 55122 52722 55134
rect 53006 55186 53058 55198
rect 53006 55122 53058 55134
rect 4734 55074 4786 55086
rect 4734 55010 4786 55022
rect 12462 55074 12514 55086
rect 12462 55010 12514 55022
rect 12910 55074 12962 55086
rect 12910 55010 12962 55022
rect 13918 55074 13970 55086
rect 13918 55010 13970 55022
rect 14702 55074 14754 55086
rect 14702 55010 14754 55022
rect 17166 55074 17218 55086
rect 17166 55010 17218 55022
rect 17502 55074 17554 55086
rect 23102 55074 23154 55086
rect 18386 55022 18398 55074
rect 18450 55022 18462 55074
rect 17502 55010 17554 55022
rect 23102 55010 23154 55022
rect 27582 55074 27634 55086
rect 27582 55010 27634 55022
rect 28366 55074 28418 55086
rect 28366 55010 28418 55022
rect 29262 55074 29314 55086
rect 29262 55010 29314 55022
rect 31726 55074 31778 55086
rect 31726 55010 31778 55022
rect 33182 55074 33234 55086
rect 33182 55010 33234 55022
rect 33406 55074 33458 55086
rect 33406 55010 33458 55022
rect 37326 55074 37378 55086
rect 37326 55010 37378 55022
rect 37998 55074 38050 55086
rect 37998 55010 38050 55022
rect 38782 55074 38834 55086
rect 38782 55010 38834 55022
rect 39118 55074 39170 55086
rect 39118 55010 39170 55022
rect 42254 55074 42306 55086
rect 42254 55010 42306 55022
rect 42590 55074 42642 55086
rect 42590 55010 42642 55022
rect 47406 55074 47458 55086
rect 47406 55010 47458 55022
rect 50766 55074 50818 55086
rect 50766 55010 50818 55022
rect 1344 54906 58576 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 58576 54906
rect 1344 54820 58576 54854
rect 14926 54738 14978 54750
rect 49982 54738 50034 54750
rect 22642 54686 22654 54738
rect 22706 54686 22718 54738
rect 26226 54686 26238 54738
rect 26290 54686 26302 54738
rect 45490 54686 45502 54738
rect 45554 54686 45566 54738
rect 14926 54674 14978 54686
rect 49982 54674 50034 54686
rect 33630 54626 33682 54638
rect 43934 54626 43986 54638
rect 16818 54574 16830 54626
rect 16882 54574 16894 54626
rect 20850 54574 20862 54626
rect 20914 54574 20926 54626
rect 21186 54574 21198 54626
rect 21250 54574 21262 54626
rect 23650 54574 23662 54626
rect 23714 54574 23726 54626
rect 23986 54574 23998 54626
rect 24050 54574 24062 54626
rect 25330 54574 25342 54626
rect 25394 54574 25406 54626
rect 37650 54574 37662 54626
rect 37714 54574 37726 54626
rect 33630 54562 33682 54574
rect 43934 54562 43986 54574
rect 46958 54626 47010 54638
rect 46958 54562 47010 54574
rect 49086 54626 49138 54638
rect 49086 54562 49138 54574
rect 50766 54626 50818 54638
rect 51874 54574 51886 54626
rect 51938 54574 51950 54626
rect 50766 54562 50818 54574
rect 13694 54514 13746 54526
rect 13694 54450 13746 54462
rect 14030 54514 14082 54526
rect 24558 54514 24610 54526
rect 26910 54514 26962 54526
rect 34526 54514 34578 54526
rect 16594 54462 16606 54514
rect 16658 54462 16670 54514
rect 17714 54462 17726 54514
rect 17778 54462 17790 54514
rect 19058 54462 19070 54514
rect 19122 54462 19134 54514
rect 19730 54462 19742 54514
rect 19794 54462 19806 54514
rect 22418 54462 22430 54514
rect 22482 54462 22494 54514
rect 25218 54462 25230 54514
rect 25282 54462 25294 54514
rect 26114 54462 26126 54514
rect 26178 54462 26190 54514
rect 28130 54462 28142 54514
rect 28194 54462 28206 54514
rect 29474 54462 29486 54514
rect 29538 54462 29550 54514
rect 30930 54462 30942 54514
rect 30994 54462 31006 54514
rect 14030 54450 14082 54462
rect 24558 54450 24610 54462
rect 26910 54450 26962 54462
rect 34526 54450 34578 54462
rect 34862 54514 34914 54526
rect 39790 54514 39842 54526
rect 41806 54514 41858 54526
rect 36082 54462 36094 54514
rect 36146 54462 36158 54514
rect 36642 54462 36654 54514
rect 36706 54462 36718 54514
rect 38210 54462 38222 54514
rect 38274 54462 38286 54514
rect 39442 54462 39454 54514
rect 39506 54462 39518 54514
rect 41234 54462 41246 54514
rect 41298 54462 41310 54514
rect 34862 54450 34914 54462
rect 39790 54450 39842 54462
rect 41806 54450 41858 54462
rect 42030 54514 42082 54526
rect 43374 54514 43426 54526
rect 45166 54514 45218 54526
rect 42130 54462 42142 54514
rect 42194 54462 42206 54514
rect 42690 54462 42702 54514
rect 42754 54462 42766 54514
rect 43698 54462 43710 54514
rect 43762 54462 43774 54514
rect 42030 54450 42082 54462
rect 43374 54450 43426 54462
rect 45166 54450 45218 54462
rect 46398 54514 46450 54526
rect 46398 54450 46450 54462
rect 46846 54514 46898 54526
rect 46846 54450 46898 54462
rect 47070 54514 47122 54526
rect 47070 54450 47122 54462
rect 47630 54514 47682 54526
rect 47630 54450 47682 54462
rect 48302 54514 48354 54526
rect 48974 54514 49026 54526
rect 50654 54514 50706 54526
rect 48738 54462 48750 54514
rect 48802 54462 48814 54514
rect 49522 54462 49534 54514
rect 49586 54462 49598 54514
rect 50194 54462 50206 54514
rect 50258 54462 50270 54514
rect 48302 54450 48354 54462
rect 48974 54450 49026 54462
rect 50654 54450 50706 54462
rect 51214 54514 51266 54526
rect 51650 54462 51662 54514
rect 51714 54462 51726 54514
rect 53218 54462 53230 54514
rect 53282 54462 53294 54514
rect 54562 54462 54574 54514
rect 54626 54462 54638 54514
rect 51214 54450 51266 54462
rect 11342 54402 11394 54414
rect 11342 54338 11394 54350
rect 11902 54402 11954 54414
rect 11902 54338 11954 54350
rect 12462 54402 12514 54414
rect 12462 54338 12514 54350
rect 12910 54402 12962 54414
rect 12910 54338 12962 54350
rect 13358 54402 13410 54414
rect 13358 54338 13410 54350
rect 13582 54402 13634 54414
rect 13582 54338 13634 54350
rect 14590 54402 14642 54414
rect 14590 54338 14642 54350
rect 15486 54402 15538 54414
rect 15486 54338 15538 54350
rect 16270 54402 16322 54414
rect 35422 54402 35474 54414
rect 41918 54402 41970 54414
rect 44494 54402 44546 54414
rect 29698 54350 29710 54402
rect 29762 54350 29774 54402
rect 31490 54350 31502 54402
rect 31554 54350 31566 54402
rect 38882 54350 38894 54402
rect 38946 54350 38958 54402
rect 39554 54350 39566 54402
rect 39618 54350 39630 54402
rect 43810 54350 43822 54402
rect 43874 54350 43886 54402
rect 16270 54338 16322 54350
rect 35422 54338 35474 54350
rect 41918 54338 41970 54350
rect 44494 54338 44546 54350
rect 44942 54402 44994 54414
rect 44942 54338 44994 54350
rect 47406 54402 47458 54414
rect 47406 54338 47458 54350
rect 50990 54402 51042 54414
rect 52882 54350 52894 54402
rect 52946 54350 52958 54402
rect 50990 54338 51042 54350
rect 24222 54290 24274 54302
rect 47854 54290 47906 54302
rect 31826 54238 31838 54290
rect 31890 54238 31902 54290
rect 38994 54238 39006 54290
rect 39058 54238 39070 54290
rect 24222 54226 24274 54238
rect 47854 54226 47906 54238
rect 49870 54290 49922 54302
rect 49870 54226 49922 54238
rect 1344 54122 58576 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 58576 54122
rect 1344 54036 58576 54070
rect 19406 53954 19458 53966
rect 16370 53902 16382 53954
rect 16434 53902 16446 53954
rect 18162 53902 18174 53954
rect 18226 53902 18238 53954
rect 19406 53890 19458 53902
rect 34078 53954 34130 53966
rect 34078 53890 34130 53902
rect 34302 53954 34354 53966
rect 34302 53890 34354 53902
rect 34750 53954 34802 53966
rect 34750 53890 34802 53902
rect 40686 53954 40738 53966
rect 40686 53890 40738 53902
rect 41470 53954 41522 53966
rect 41470 53890 41522 53902
rect 42814 53954 42866 53966
rect 42814 53890 42866 53902
rect 43262 53954 43314 53966
rect 43262 53890 43314 53902
rect 12462 53842 12514 53854
rect 35198 53842 35250 53854
rect 40798 53842 40850 53854
rect 18050 53790 18062 53842
rect 18114 53790 18126 53842
rect 20402 53790 20414 53842
rect 20466 53790 20478 53842
rect 35410 53790 35422 53842
rect 35474 53790 35486 53842
rect 40002 53790 40014 53842
rect 40066 53790 40078 53842
rect 12462 53778 12514 53790
rect 35198 53778 35250 53790
rect 40798 53778 40850 53790
rect 9998 53730 10050 53742
rect 9538 53678 9550 53730
rect 9602 53678 9614 53730
rect 9998 53666 10050 53678
rect 12798 53730 12850 53742
rect 12798 53666 12850 53678
rect 13918 53730 13970 53742
rect 13918 53666 13970 53678
rect 14478 53730 14530 53742
rect 14478 53666 14530 53678
rect 15374 53730 15426 53742
rect 15374 53666 15426 53678
rect 15710 53730 15762 53742
rect 19630 53730 19682 53742
rect 30158 53730 30210 53742
rect 33854 53730 33906 53742
rect 36878 53730 36930 53742
rect 15922 53678 15934 53730
rect 15986 53678 15998 53730
rect 16930 53678 16942 53730
rect 16994 53678 17006 53730
rect 20514 53678 20526 53730
rect 20578 53678 20590 53730
rect 21522 53678 21534 53730
rect 21586 53678 21598 53730
rect 24098 53678 24110 53730
rect 24162 53678 24174 53730
rect 26450 53678 26462 53730
rect 26514 53678 26526 53730
rect 26674 53678 26686 53730
rect 26738 53678 26750 53730
rect 27682 53678 27694 53730
rect 27746 53678 27758 53730
rect 28354 53678 28366 53730
rect 28418 53678 28430 53730
rect 30594 53678 30606 53730
rect 30658 53678 30670 53730
rect 32274 53678 32286 53730
rect 32338 53678 32350 53730
rect 33058 53678 33070 53730
rect 33122 53678 33134 53730
rect 35522 53678 35534 53730
rect 35586 53678 35598 53730
rect 15710 53666 15762 53678
rect 19630 53666 19682 53678
rect 30158 53666 30210 53678
rect 33854 53666 33906 53678
rect 36878 53666 36930 53678
rect 37214 53730 37266 53742
rect 42254 53730 42306 53742
rect 39666 53678 39678 53730
rect 39730 53678 39742 53730
rect 37214 53666 37266 53678
rect 42254 53666 42306 53678
rect 42478 53730 42530 53742
rect 42478 53666 42530 53678
rect 47182 53730 47234 53742
rect 47182 53666 47234 53678
rect 47742 53730 47794 53742
rect 47742 53666 47794 53678
rect 47966 53730 48018 53742
rect 55570 53678 55582 53730
rect 55634 53678 55646 53730
rect 47966 53666 48018 53678
rect 17390 53618 17442 53630
rect 29150 53618 29202 53630
rect 11890 53566 11902 53618
rect 11954 53566 11966 53618
rect 12226 53566 12238 53618
rect 12290 53566 12302 53618
rect 17826 53566 17838 53618
rect 17890 53566 17902 53618
rect 22418 53566 22430 53618
rect 22482 53566 22494 53618
rect 23426 53566 23438 53618
rect 23490 53566 23502 53618
rect 28578 53566 28590 53618
rect 28642 53566 28654 53618
rect 17390 53554 17442 53566
rect 29150 53554 29202 53566
rect 29822 53618 29874 53630
rect 29822 53554 29874 53566
rect 29934 53618 29986 53630
rect 37550 53618 37602 53630
rect 31602 53566 31614 53618
rect 31666 53566 31678 53618
rect 32162 53566 32174 53618
rect 32226 53566 32238 53618
rect 29934 53554 29986 53566
rect 37550 53554 37602 53566
rect 37998 53618 38050 53630
rect 37998 53554 38050 53566
rect 40350 53618 40402 53630
rect 40350 53554 40402 53566
rect 41358 53618 41410 53630
rect 41358 53554 41410 53566
rect 43150 53618 43202 53630
rect 43150 53554 43202 53566
rect 43262 53618 43314 53630
rect 43262 53554 43314 53566
rect 47630 53618 47682 53630
rect 47630 53554 47682 53566
rect 49086 53618 49138 53630
rect 49086 53554 49138 53566
rect 50990 53618 51042 53630
rect 50990 53554 51042 53566
rect 53566 53618 53618 53630
rect 53566 53554 53618 53566
rect 53902 53618 53954 53630
rect 57250 53566 57262 53618
rect 57314 53566 57326 53618
rect 53902 53554 53954 53566
rect 10894 53506 10946 53518
rect 10894 53442 10946 53454
rect 11342 53506 11394 53518
rect 11342 53442 11394 53454
rect 13694 53506 13746 53518
rect 13694 53442 13746 53454
rect 14814 53506 14866 53518
rect 14814 53442 14866 53454
rect 20638 53506 20690 53518
rect 27358 53506 27410 53518
rect 35982 53506 36034 53518
rect 24322 53454 24334 53506
rect 24386 53454 24398 53506
rect 28018 53454 28030 53506
rect 28082 53454 28094 53506
rect 29474 53454 29486 53506
rect 29538 53454 29550 53506
rect 31714 53454 31726 53506
rect 31778 53454 31790 53506
rect 33170 53454 33182 53506
rect 33234 53454 33246 53506
rect 20638 53442 20690 53454
rect 27358 53442 27410 53454
rect 35982 53442 36034 53454
rect 36430 53506 36482 53518
rect 36430 53442 36482 53454
rect 37214 53506 37266 53518
rect 37214 53442 37266 53454
rect 39006 53506 39058 53518
rect 39006 53442 39058 53454
rect 40910 53506 40962 53518
rect 40910 53442 40962 53454
rect 41470 53506 41522 53518
rect 41470 53442 41522 53454
rect 51102 53506 51154 53518
rect 51102 53442 51154 53454
rect 51326 53506 51378 53518
rect 51326 53442 51378 53454
rect 1344 53338 58576 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 58576 53338
rect 1344 53252 58576 53286
rect 13358 53170 13410 53182
rect 13358 53106 13410 53118
rect 17502 53170 17554 53182
rect 17502 53106 17554 53118
rect 18846 53170 18898 53182
rect 18846 53106 18898 53118
rect 22766 53170 22818 53182
rect 22766 53106 22818 53118
rect 24334 53170 24386 53182
rect 24334 53106 24386 53118
rect 26014 53170 26066 53182
rect 26014 53106 26066 53118
rect 31950 53170 32002 53182
rect 33630 53170 33682 53182
rect 32274 53118 32286 53170
rect 32338 53118 32350 53170
rect 31950 53106 32002 53118
rect 33630 53106 33682 53118
rect 34078 53170 34130 53182
rect 34078 53106 34130 53118
rect 35422 53170 35474 53182
rect 35422 53106 35474 53118
rect 37998 53170 38050 53182
rect 37998 53106 38050 53118
rect 38894 53170 38946 53182
rect 38894 53106 38946 53118
rect 39566 53170 39618 53182
rect 39566 53106 39618 53118
rect 39790 53170 39842 53182
rect 39790 53106 39842 53118
rect 40126 53170 40178 53182
rect 50866 53118 50878 53170
rect 50930 53118 50942 53170
rect 40126 53106 40178 53118
rect 23550 53058 23602 53070
rect 34974 53058 35026 53070
rect 22530 53006 22542 53058
rect 22594 53006 22606 53058
rect 23202 53006 23214 53058
rect 23266 53006 23278 53058
rect 24658 53006 24670 53058
rect 24722 53006 24734 53058
rect 27906 53006 27918 53058
rect 27970 53006 27982 53058
rect 23550 52994 23602 53006
rect 34974 52994 35026 53006
rect 39454 53058 39506 53070
rect 39454 52994 39506 53006
rect 46510 53058 46562 53070
rect 53454 53058 53506 53070
rect 51538 53006 51550 53058
rect 51602 53006 51614 53058
rect 46510 52994 46562 53006
rect 53454 52994 53506 53006
rect 12574 52946 12626 52958
rect 18510 52946 18562 52958
rect 50318 52946 50370 52958
rect 10322 52894 10334 52946
rect 10386 52894 10398 52946
rect 12114 52894 12126 52946
rect 12178 52894 12190 52946
rect 14242 52894 14254 52946
rect 14306 52894 14318 52946
rect 15922 52894 15934 52946
rect 15986 52894 15998 52946
rect 19170 52894 19182 52946
rect 19234 52894 19246 52946
rect 19730 52894 19742 52946
rect 19794 52894 19806 52946
rect 21298 52894 21310 52946
rect 21362 52894 21374 52946
rect 28466 52894 28478 52946
rect 28530 52894 28542 52946
rect 29474 52894 29486 52946
rect 29538 52894 29550 52946
rect 30706 52894 30718 52946
rect 30770 52894 30782 52946
rect 45938 52894 45950 52946
rect 46002 52894 46014 52946
rect 50082 52894 50094 52946
rect 50146 52894 50158 52946
rect 12574 52882 12626 52894
rect 18510 52882 18562 52894
rect 50318 52882 50370 52894
rect 50430 52946 50482 52958
rect 52770 52894 52782 52946
rect 52834 52894 52846 52946
rect 50430 52882 50482 52894
rect 13806 52834 13858 52846
rect 18062 52834 18114 52846
rect 11442 52782 11454 52834
rect 11506 52782 11518 52834
rect 14130 52782 14142 52834
rect 14194 52782 14206 52834
rect 16370 52782 16382 52834
rect 16434 52782 16446 52834
rect 13806 52770 13858 52782
rect 18062 52770 18114 52782
rect 24110 52834 24162 52846
rect 24110 52770 24162 52782
rect 25566 52834 25618 52846
rect 25566 52770 25618 52782
rect 26574 52834 26626 52846
rect 26574 52770 26626 52782
rect 27022 52834 27074 52846
rect 33182 52834 33234 52846
rect 28914 52782 28926 52834
rect 28978 52782 28990 52834
rect 27022 52770 27074 52782
rect 33182 52770 33234 52782
rect 34526 52834 34578 52846
rect 34526 52770 34578 52782
rect 38446 52834 38498 52846
rect 38446 52770 38498 52782
rect 41806 52834 41858 52846
rect 45714 52782 45726 52834
rect 45778 52782 45790 52834
rect 51314 52782 51326 52834
rect 51378 52782 51390 52834
rect 41806 52770 41858 52782
rect 32946 52670 32958 52722
rect 33010 52719 33022 52722
rect 33506 52719 33518 52722
rect 33010 52673 33518 52719
rect 33010 52670 33022 52673
rect 33506 52670 33518 52673
rect 33570 52670 33582 52722
rect 33842 52670 33854 52722
rect 33906 52719 33918 52722
rect 34626 52719 34638 52722
rect 33906 52673 34638 52719
rect 33906 52670 33918 52673
rect 34626 52670 34638 52673
rect 34690 52670 34702 52722
rect 1344 52554 58576 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 58576 52554
rect 1344 52468 58576 52502
rect 19406 52386 19458 52398
rect 45838 52386 45890 52398
rect 11106 52334 11118 52386
rect 11170 52334 11182 52386
rect 13458 52334 13470 52386
rect 13522 52383 13534 52386
rect 13794 52383 13806 52386
rect 13522 52337 13806 52383
rect 13522 52334 13534 52337
rect 13794 52334 13806 52337
rect 13858 52334 13870 52386
rect 28018 52334 28030 52386
rect 28082 52334 28094 52386
rect 35746 52334 35758 52386
rect 35810 52334 35822 52386
rect 41682 52334 41694 52386
rect 41746 52334 41758 52386
rect 19406 52322 19458 52334
rect 45838 52322 45890 52334
rect 8094 52274 8146 52286
rect 9774 52274 9826 52286
rect 13806 52274 13858 52286
rect 18286 52274 18338 52286
rect 8754 52222 8766 52274
rect 8818 52222 8830 52274
rect 10658 52222 10670 52274
rect 10722 52222 10734 52274
rect 12338 52222 12350 52274
rect 12402 52222 12414 52274
rect 17602 52222 17614 52274
rect 17666 52222 17678 52274
rect 8094 52210 8146 52222
rect 9774 52210 9826 52222
rect 13806 52210 13858 52222
rect 18286 52210 18338 52222
rect 23326 52274 23378 52286
rect 23326 52210 23378 52222
rect 23774 52274 23826 52286
rect 29598 52274 29650 52286
rect 27570 52222 27582 52274
rect 27634 52222 27646 52274
rect 23774 52210 23826 52222
rect 29598 52210 29650 52222
rect 31838 52274 31890 52286
rect 38558 52274 38610 52286
rect 33842 52222 33854 52274
rect 33906 52222 33918 52274
rect 37426 52222 37438 52274
rect 37490 52222 37502 52274
rect 31838 52210 31890 52222
rect 38558 52210 38610 52222
rect 39006 52274 39058 52286
rect 39006 52210 39058 52222
rect 43262 52274 43314 52286
rect 43262 52210 43314 52222
rect 44046 52274 44098 52286
rect 44046 52210 44098 52222
rect 45278 52274 45330 52286
rect 45278 52210 45330 52222
rect 48190 52274 48242 52286
rect 48190 52210 48242 52222
rect 8318 52162 8370 52174
rect 18622 52162 18674 52174
rect 9314 52110 9326 52162
rect 9378 52110 9390 52162
rect 10434 52110 10446 52162
rect 10498 52110 10510 52162
rect 10770 52110 10782 52162
rect 10834 52110 10846 52162
rect 12562 52110 12574 52162
rect 12626 52110 12638 52162
rect 14354 52110 14366 52162
rect 14418 52110 14430 52162
rect 15810 52110 15822 52162
rect 15874 52110 15886 52162
rect 16146 52110 16158 52162
rect 16210 52110 16222 52162
rect 8318 52098 8370 52110
rect 18622 52098 18674 52110
rect 20302 52162 20354 52174
rect 20302 52098 20354 52110
rect 20414 52162 20466 52174
rect 20414 52098 20466 52110
rect 20750 52162 20802 52174
rect 29038 52162 29090 52174
rect 21410 52110 21422 52162
rect 21474 52110 21486 52162
rect 22530 52110 22542 52162
rect 22594 52110 22606 52162
rect 24210 52110 24222 52162
rect 24274 52110 24286 52162
rect 24434 52110 24446 52162
rect 24498 52110 24510 52162
rect 26002 52110 26014 52162
rect 26066 52110 26078 52162
rect 27122 52110 27134 52162
rect 27186 52110 27198 52162
rect 20750 52098 20802 52110
rect 29038 52098 29090 52110
rect 30606 52162 30658 52174
rect 32734 52162 32786 52174
rect 30818 52110 30830 52162
rect 30882 52110 30894 52162
rect 31154 52110 31166 52162
rect 31218 52110 31230 52162
rect 32162 52110 32174 52162
rect 32226 52110 32238 52162
rect 30606 52098 30658 52110
rect 32734 52098 32786 52110
rect 33406 52162 33458 52174
rect 33406 52098 33458 52110
rect 34302 52162 34354 52174
rect 34302 52098 34354 52110
rect 34526 52162 34578 52174
rect 34526 52098 34578 52110
rect 35198 52162 35250 52174
rect 35198 52098 35250 52110
rect 35422 52162 35474 52174
rect 41022 52162 41074 52174
rect 37202 52110 37214 52162
rect 37266 52110 37278 52162
rect 39442 52110 39454 52162
rect 39506 52110 39518 52162
rect 40002 52110 40014 52162
rect 40066 52110 40078 52162
rect 35422 52098 35474 52110
rect 41022 52098 41074 52110
rect 41134 52162 41186 52174
rect 41134 52098 41186 52110
rect 41246 52162 41298 52174
rect 41246 52098 41298 52110
rect 43598 52162 43650 52174
rect 43598 52098 43650 52110
rect 43822 52162 43874 52174
rect 43822 52098 43874 52110
rect 44830 52162 44882 52174
rect 44830 52098 44882 52110
rect 45726 52162 45778 52174
rect 50978 52110 50990 52162
rect 51042 52110 51054 52162
rect 51874 52110 51886 52162
rect 51938 52110 51950 52162
rect 45726 52098 45778 52110
rect 38110 52050 38162 52062
rect 43486 52050 43538 52062
rect 12450 51998 12462 52050
rect 12514 51998 12526 52050
rect 17154 51998 17166 52050
rect 17218 51998 17230 52050
rect 21522 51998 21534 52050
rect 21586 51998 21598 52050
rect 40114 51998 40126 52050
rect 40178 51998 40190 52050
rect 38110 51986 38162 51998
rect 43486 51986 43538 51998
rect 45054 52050 45106 52062
rect 45054 51986 45106 51998
rect 45390 52050 45442 52062
rect 51202 51998 51214 52050
rect 51266 51998 51278 52050
rect 45390 51986 45442 51998
rect 20638 51938 20690 51950
rect 29486 51938 29538 51950
rect 22306 51886 22318 51938
rect 22370 51886 22382 51938
rect 20638 51874 20690 51886
rect 29486 51874 29538 51886
rect 29710 51938 29762 51950
rect 29710 51874 29762 51886
rect 30382 51938 30434 51950
rect 38446 51938 38498 51950
rect 45838 51938 45890 51950
rect 34850 51886 34862 51938
rect 34914 51886 34926 51938
rect 39666 51886 39678 51938
rect 39730 51886 39742 51938
rect 30382 51874 30434 51886
rect 38446 51874 38498 51886
rect 45838 51874 45890 51886
rect 46734 51938 46786 51950
rect 46734 51874 46786 51886
rect 47182 51938 47234 51950
rect 47182 51874 47234 51886
rect 47630 51938 47682 51950
rect 51986 51886 51998 51938
rect 52050 51886 52062 51938
rect 47630 51874 47682 51886
rect 1344 51770 58576 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 58576 51770
rect 1344 51684 58576 51718
rect 22990 51602 23042 51614
rect 21858 51550 21870 51602
rect 21922 51550 21934 51602
rect 22990 51538 23042 51550
rect 25230 51602 25282 51614
rect 25230 51538 25282 51550
rect 31166 51602 31218 51614
rect 39902 51602 39954 51614
rect 31714 51550 31726 51602
rect 31778 51550 31790 51602
rect 31166 51538 31218 51550
rect 39902 51538 39954 51550
rect 40126 51602 40178 51614
rect 44034 51550 44046 51602
rect 44098 51550 44110 51602
rect 40126 51538 40178 51550
rect 1710 51490 1762 51502
rect 1710 51426 1762 51438
rect 9998 51490 10050 51502
rect 9998 51426 10050 51438
rect 13918 51490 13970 51502
rect 13918 51426 13970 51438
rect 25678 51490 25730 51502
rect 29822 51490 29874 51502
rect 38446 51490 38498 51502
rect 26898 51438 26910 51490
rect 26962 51438 26974 51490
rect 34850 51438 34862 51490
rect 34914 51438 34926 51490
rect 35298 51438 35310 51490
rect 35362 51438 35374 51490
rect 25678 51426 25730 51438
rect 29822 51426 29874 51438
rect 38446 51426 38498 51438
rect 39678 51490 39730 51502
rect 39678 51426 39730 51438
rect 42702 51490 42754 51502
rect 42702 51426 42754 51438
rect 43038 51490 43090 51502
rect 55022 51490 55074 51502
rect 46162 51438 46174 51490
rect 46226 51438 46238 51490
rect 50418 51438 50430 51490
rect 50482 51438 50494 51490
rect 43038 51426 43090 51438
rect 55022 51426 55074 51438
rect 12686 51378 12738 51390
rect 10322 51326 10334 51378
rect 10386 51326 10398 51378
rect 11106 51326 11118 51378
rect 11170 51326 11182 51378
rect 12686 51314 12738 51326
rect 15486 51378 15538 51390
rect 20078 51378 20130 51390
rect 16370 51326 16382 51378
rect 16434 51326 16446 51378
rect 17714 51326 17726 51378
rect 17778 51326 17790 51378
rect 18834 51326 18846 51378
rect 18898 51326 18910 51378
rect 19170 51326 19182 51378
rect 19234 51326 19246 51378
rect 19618 51326 19630 51378
rect 19682 51326 19694 51378
rect 15486 51314 15538 51326
rect 20078 51314 20130 51326
rect 20638 51378 20690 51390
rect 20638 51314 20690 51326
rect 20750 51378 20802 51390
rect 20750 51314 20802 51326
rect 20862 51378 20914 51390
rect 21534 51378 21586 51390
rect 22878 51378 22930 51390
rect 30942 51378 30994 51390
rect 21186 51326 21198 51378
rect 21250 51326 21262 51378
rect 22530 51326 22542 51378
rect 22594 51326 22606 51378
rect 24210 51326 24222 51378
rect 24274 51326 24286 51378
rect 25442 51326 25454 51378
rect 25506 51326 25518 51378
rect 26114 51326 26126 51378
rect 26178 51326 26190 51378
rect 27122 51326 27134 51378
rect 27186 51326 27198 51378
rect 28690 51326 28702 51378
rect 28754 51326 28766 51378
rect 29026 51326 29038 51378
rect 29090 51326 29102 51378
rect 30706 51326 30718 51378
rect 30770 51326 30782 51378
rect 20862 51314 20914 51326
rect 21534 51314 21586 51326
rect 22878 51314 22930 51326
rect 30942 51314 30994 51326
rect 31278 51378 31330 51390
rect 36878 51378 36930 51390
rect 33730 51326 33742 51378
rect 33794 51326 33806 51378
rect 34178 51326 34190 51378
rect 34242 51326 34254 51378
rect 31278 51314 31330 51326
rect 36878 51314 36930 51326
rect 37326 51378 37378 51390
rect 37326 51314 37378 51326
rect 40350 51378 40402 51390
rect 48638 51378 48690 51390
rect 47506 51326 47518 51378
rect 47570 51326 47582 51378
rect 40350 51314 40402 51326
rect 48638 51314 48690 51326
rect 49198 51378 49250 51390
rect 49198 51314 49250 51326
rect 49422 51378 49474 51390
rect 49422 51314 49474 51326
rect 54686 51378 54738 51390
rect 54686 51314 54738 51326
rect 23886 51266 23938 51278
rect 26574 51266 26626 51278
rect 32286 51266 32338 51278
rect 10658 51214 10670 51266
rect 10722 51214 10734 51266
rect 12226 51214 12238 51266
rect 12290 51214 12302 51266
rect 13234 51214 13246 51266
rect 13298 51214 13310 51266
rect 14242 51214 14254 51266
rect 14306 51214 14318 51266
rect 16706 51214 16718 51266
rect 16770 51214 16782 51266
rect 17826 51214 17838 51266
rect 17890 51214 17902 51266
rect 24546 51214 24558 51266
rect 24610 51214 24622 51266
rect 31154 51214 31166 51266
rect 31218 51214 31230 51266
rect 23886 51202 23938 51214
rect 26574 51202 26626 51214
rect 32286 51202 32338 51214
rect 33182 51266 33234 51278
rect 43486 51266 43538 51278
rect 34514 51214 34526 51266
rect 34578 51214 34590 51266
rect 36530 51214 36542 51266
rect 36594 51214 36606 51266
rect 33182 51202 33234 51214
rect 43486 51202 43538 51214
rect 46510 51266 46562 51278
rect 46510 51202 46562 51214
rect 46958 51266 47010 51278
rect 46958 51202 47010 51214
rect 47966 51266 48018 51278
rect 47966 51202 48018 51214
rect 15598 51154 15650 51166
rect 14466 51102 14478 51154
rect 14530 51102 14542 51154
rect 15598 51090 15650 51102
rect 18622 51154 18674 51166
rect 22206 51154 22258 51166
rect 20066 51102 20078 51154
rect 20130 51102 20142 51154
rect 18622 51090 18674 51102
rect 22206 51090 22258 51102
rect 22542 51154 22594 51166
rect 22542 51090 22594 51102
rect 22990 51154 23042 51166
rect 22990 51090 23042 51102
rect 25566 51154 25618 51166
rect 25566 51090 25618 51102
rect 32062 51154 32114 51166
rect 32062 51090 32114 51102
rect 40238 51154 40290 51166
rect 40238 51090 40290 51102
rect 43710 51154 43762 51166
rect 43710 51090 43762 51102
rect 48862 51154 48914 51166
rect 48862 51090 48914 51102
rect 1344 50986 58576 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 58576 50986
rect 1344 50900 58576 50934
rect 28366 50818 28418 50830
rect 14130 50766 14142 50818
rect 14194 50766 14206 50818
rect 24994 50766 25006 50818
rect 25058 50766 25070 50818
rect 28366 50754 28418 50766
rect 29822 50818 29874 50830
rect 29822 50754 29874 50766
rect 30158 50818 30210 50830
rect 30158 50754 30210 50766
rect 31726 50818 31778 50830
rect 31726 50754 31778 50766
rect 32958 50818 33010 50830
rect 32958 50754 33010 50766
rect 37550 50818 37602 50830
rect 37550 50754 37602 50766
rect 37998 50818 38050 50830
rect 37998 50754 38050 50766
rect 38110 50818 38162 50830
rect 38110 50754 38162 50766
rect 48638 50818 48690 50830
rect 48638 50754 48690 50766
rect 52894 50818 52946 50830
rect 52894 50754 52946 50766
rect 9550 50706 9602 50718
rect 9550 50642 9602 50654
rect 12462 50706 12514 50718
rect 16718 50706 16770 50718
rect 29486 50706 29538 50718
rect 13570 50654 13582 50706
rect 13634 50654 13646 50706
rect 15026 50654 15038 50706
rect 15090 50654 15102 50706
rect 24882 50654 24894 50706
rect 24946 50654 24958 50706
rect 12462 50642 12514 50654
rect 16718 50642 16770 50654
rect 29486 50642 29538 50654
rect 30942 50706 30994 50718
rect 30942 50642 30994 50654
rect 33294 50706 33346 50718
rect 33294 50642 33346 50654
rect 39230 50706 39282 50718
rect 39230 50642 39282 50654
rect 39678 50706 39730 50718
rect 52670 50706 52722 50718
rect 43698 50654 43710 50706
rect 43762 50654 43774 50706
rect 49634 50654 49646 50706
rect 49698 50654 49710 50706
rect 39678 50642 39730 50654
rect 52670 50642 52722 50654
rect 53230 50706 53282 50718
rect 54574 50706 54626 50718
rect 53666 50654 53678 50706
rect 53730 50654 53742 50706
rect 53230 50642 53282 50654
rect 54574 50642 54626 50654
rect 57934 50706 57986 50718
rect 57934 50642 57986 50654
rect 16046 50594 16098 50606
rect 9090 50542 9102 50594
rect 9154 50542 9166 50594
rect 13682 50542 13694 50594
rect 13746 50542 13758 50594
rect 15586 50542 15598 50594
rect 15650 50542 15662 50594
rect 16046 50530 16098 50542
rect 16942 50594 16994 50606
rect 16942 50530 16994 50542
rect 17502 50594 17554 50606
rect 19630 50594 19682 50606
rect 28030 50594 28082 50606
rect 18386 50542 18398 50594
rect 18450 50542 18462 50594
rect 18722 50542 18734 50594
rect 18786 50542 18798 50594
rect 20290 50542 20302 50594
rect 20354 50542 20366 50594
rect 21298 50542 21310 50594
rect 21362 50542 21374 50594
rect 21634 50542 21646 50594
rect 21698 50542 21710 50594
rect 23650 50542 23662 50594
rect 23714 50542 23726 50594
rect 24322 50542 24334 50594
rect 24386 50542 24398 50594
rect 27346 50542 27358 50594
rect 27410 50542 27422 50594
rect 17502 50530 17554 50542
rect 19630 50530 19682 50542
rect 28030 50530 28082 50542
rect 30830 50594 30882 50606
rect 30830 50530 30882 50542
rect 31054 50594 31106 50606
rect 31054 50530 31106 50542
rect 32286 50594 32338 50606
rect 32286 50530 32338 50542
rect 33742 50594 33794 50606
rect 33742 50530 33794 50542
rect 36318 50594 36370 50606
rect 36318 50530 36370 50542
rect 37326 50594 37378 50606
rect 37326 50530 37378 50542
rect 37998 50594 38050 50606
rect 37998 50530 38050 50542
rect 42478 50594 42530 50606
rect 45614 50594 45666 50606
rect 43362 50542 43374 50594
rect 43426 50542 43438 50594
rect 42478 50530 42530 50542
rect 45614 50530 45666 50542
rect 46174 50594 46226 50606
rect 48862 50594 48914 50606
rect 46498 50542 46510 50594
rect 46562 50542 46574 50594
rect 47282 50542 47294 50594
rect 47346 50542 47358 50594
rect 46174 50530 46226 50542
rect 48862 50530 48914 50542
rect 49086 50594 49138 50606
rect 49086 50530 49138 50542
rect 50094 50594 50146 50606
rect 50094 50530 50146 50542
rect 50654 50594 50706 50606
rect 53890 50542 53902 50594
rect 53954 50542 53966 50594
rect 55570 50542 55582 50594
rect 55634 50542 55646 50594
rect 50654 50530 50706 50542
rect 19742 50482 19794 50494
rect 8194 50430 8206 50482
rect 8258 50430 8270 50482
rect 17826 50430 17838 50482
rect 17890 50430 17902 50482
rect 19742 50418 19794 50430
rect 20750 50482 20802 50494
rect 20750 50418 20802 50430
rect 26462 50482 26514 50494
rect 30046 50482 30098 50494
rect 27458 50430 27470 50482
rect 27522 50430 27534 50482
rect 26462 50418 26514 50430
rect 30046 50418 30098 50430
rect 31390 50482 31442 50494
rect 31390 50418 31442 50430
rect 31614 50482 31666 50494
rect 31614 50418 31666 50430
rect 32846 50482 32898 50494
rect 32846 50418 32898 50430
rect 35758 50482 35810 50494
rect 35758 50418 35810 50430
rect 42142 50482 42194 50494
rect 42142 50418 42194 50430
rect 44270 50482 44322 50494
rect 44270 50418 44322 50430
rect 46734 50482 46786 50494
rect 46734 50418 46786 50430
rect 46846 50482 46898 50494
rect 46846 50418 46898 50430
rect 48078 50482 48130 50494
rect 48078 50418 48130 50430
rect 48414 50482 48466 50494
rect 48414 50418 48466 50430
rect 50206 50482 50258 50494
rect 50206 50418 50258 50430
rect 50766 50482 50818 50494
rect 50766 50418 50818 50430
rect 54910 50482 54962 50494
rect 54910 50418 54962 50430
rect 55246 50482 55298 50494
rect 55246 50418 55298 50430
rect 7870 50370 7922 50382
rect 7870 50306 7922 50318
rect 8766 50370 8818 50382
rect 8766 50306 8818 50318
rect 10334 50370 10386 50382
rect 10334 50306 10386 50318
rect 10782 50370 10834 50382
rect 10782 50306 10834 50318
rect 11118 50370 11170 50382
rect 11118 50306 11170 50318
rect 11678 50370 11730 50382
rect 11678 50306 11730 50318
rect 12014 50370 12066 50382
rect 12014 50306 12066 50318
rect 13022 50370 13074 50382
rect 13022 50306 13074 50318
rect 14590 50370 14642 50382
rect 19966 50370 20018 50382
rect 18722 50318 18734 50370
rect 18786 50318 18798 50370
rect 14590 50306 14642 50318
rect 19966 50306 20018 50318
rect 26910 50370 26962 50382
rect 26910 50306 26962 50318
rect 30606 50370 30658 50382
rect 30606 50306 30658 50318
rect 32622 50370 32674 50382
rect 50990 50370 51042 50382
rect 42802 50318 42814 50370
rect 42866 50318 42878 50370
rect 32622 50306 32674 50318
rect 50990 50306 51042 50318
rect 1344 50202 58576 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 58576 50202
rect 1344 50116 58576 50150
rect 15262 50034 15314 50046
rect 8530 49982 8542 50034
rect 8594 49982 8606 50034
rect 15262 49970 15314 49982
rect 16830 50034 16882 50046
rect 31614 50034 31666 50046
rect 22866 49982 22878 50034
rect 22930 49982 22942 50034
rect 29698 49982 29710 50034
rect 29762 49982 29774 50034
rect 16830 49970 16882 49982
rect 31614 49970 31666 49982
rect 33630 50034 33682 50046
rect 33630 49970 33682 49982
rect 36094 50034 36146 50046
rect 36094 49970 36146 49982
rect 41022 50034 41074 50046
rect 41022 49970 41074 49982
rect 41470 50034 41522 50046
rect 46946 49982 46958 50034
rect 47010 49982 47022 50034
rect 41470 49970 41522 49982
rect 13358 49922 13410 49934
rect 31278 49922 31330 49934
rect 18722 49870 18734 49922
rect 18786 49870 18798 49922
rect 20178 49870 20190 49922
rect 20242 49870 20254 49922
rect 21410 49870 21422 49922
rect 21474 49870 21486 49922
rect 23650 49870 23662 49922
rect 23714 49870 23726 49922
rect 24658 49870 24670 49922
rect 24722 49870 24734 49922
rect 26562 49870 26574 49922
rect 26626 49870 26638 49922
rect 30370 49870 30382 49922
rect 30434 49870 30446 49922
rect 13358 49858 13410 49870
rect 31278 49858 31330 49870
rect 31502 49922 31554 49934
rect 31502 49858 31554 49870
rect 32398 49922 32450 49934
rect 54910 49922 54962 49934
rect 35186 49870 35198 49922
rect 35250 49870 35262 49922
rect 43474 49870 43486 49922
rect 43538 49870 43550 49922
rect 44370 49870 44382 49922
rect 44434 49870 44446 49922
rect 46162 49870 46174 49922
rect 46226 49870 46238 49922
rect 50978 49870 50990 49922
rect 51042 49870 51054 49922
rect 52322 49870 52334 49922
rect 52386 49870 52398 49922
rect 32398 49858 32450 49870
rect 54910 49858 54962 49870
rect 8878 49810 8930 49822
rect 8306 49758 8318 49810
rect 8370 49758 8382 49810
rect 8878 49746 8930 49758
rect 9550 49810 9602 49822
rect 11342 49810 11394 49822
rect 14142 49810 14194 49822
rect 24334 49810 24386 49822
rect 31726 49810 31778 49822
rect 10994 49758 11006 49810
rect 11058 49758 11070 49810
rect 12338 49758 12350 49810
rect 12402 49758 12414 49810
rect 17378 49758 17390 49810
rect 17442 49758 17454 49810
rect 17938 49758 17950 49810
rect 18002 49758 18014 49810
rect 18498 49758 18510 49810
rect 18562 49758 18574 49810
rect 19282 49758 19294 49810
rect 19346 49758 19358 49810
rect 19842 49758 19854 49810
rect 19906 49758 19918 49810
rect 21634 49758 21646 49810
rect 21698 49758 21710 49810
rect 22754 49758 22766 49810
rect 22818 49758 22830 49810
rect 25442 49758 25454 49810
rect 25506 49758 25518 49810
rect 27234 49758 27246 49810
rect 27298 49758 27310 49810
rect 27794 49758 27806 49810
rect 27858 49758 27870 49810
rect 29362 49758 29374 49810
rect 29426 49758 29438 49810
rect 9550 49746 9602 49758
rect 11342 49746 11394 49758
rect 14142 49746 14194 49758
rect 24334 49746 24386 49758
rect 31726 49746 31778 49758
rect 31838 49810 31890 49822
rect 31838 49746 31890 49758
rect 33518 49810 33570 49822
rect 33518 49746 33570 49758
rect 33854 49810 33906 49822
rect 36654 49810 36706 49822
rect 40238 49810 40290 49822
rect 34290 49758 34302 49810
rect 34354 49758 34366 49810
rect 35410 49758 35422 49810
rect 35474 49758 35486 49810
rect 39330 49758 39342 49810
rect 39394 49758 39406 49810
rect 33854 49746 33906 49758
rect 36654 49746 36706 49758
rect 40238 49746 40290 49758
rect 42142 49810 42194 49822
rect 51774 49810 51826 49822
rect 45266 49758 45278 49810
rect 45330 49758 45342 49810
rect 45938 49758 45950 49810
rect 46002 49758 46014 49810
rect 46834 49758 46846 49810
rect 46898 49758 46910 49810
rect 42142 49746 42194 49758
rect 51774 49746 51826 49758
rect 53902 49810 53954 49822
rect 53902 49746 53954 49758
rect 54350 49810 54402 49822
rect 54350 49746 54402 49758
rect 8990 49698 9042 49710
rect 11454 49698 11506 49710
rect 9986 49646 9998 49698
rect 10050 49646 10062 49698
rect 8990 49634 9042 49646
rect 11454 49634 11506 49646
rect 12014 49698 12066 49710
rect 12014 49634 12066 49646
rect 14702 49698 14754 49710
rect 14702 49634 14754 49646
rect 15822 49698 15874 49710
rect 15822 49634 15874 49646
rect 16382 49698 16434 49710
rect 16382 49634 16434 49646
rect 18286 49698 18338 49710
rect 37998 49698 38050 49710
rect 19954 49646 19966 49698
rect 20018 49646 20030 49698
rect 34290 49695 34302 49698
rect 33969 49649 34302 49695
rect 18286 49634 18338 49646
rect 33969 49586 34015 49649
rect 34290 49646 34302 49649
rect 34354 49646 34366 49698
rect 34962 49646 34974 49698
rect 35026 49646 35038 49698
rect 39778 49646 39790 49698
rect 39842 49646 39854 49698
rect 50866 49646 50878 49698
rect 50930 49646 50942 49698
rect 54002 49646 54014 49698
rect 54066 49646 54078 49698
rect 37998 49634 38050 49646
rect 45166 49586 45218 49598
rect 33954 49534 33966 49586
rect 34018 49534 34030 49586
rect 45166 49522 45218 49534
rect 1344 49418 58576 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 58576 49418
rect 1344 49332 58576 49366
rect 9886 49250 9938 49262
rect 33506 49247 33518 49250
rect 9886 49186 9938 49198
rect 33073 49201 33518 49247
rect 1934 49138 1986 49150
rect 1934 49074 1986 49086
rect 10558 49138 10610 49150
rect 10558 49074 10610 49086
rect 11006 49138 11058 49150
rect 20190 49138 20242 49150
rect 24222 49138 24274 49150
rect 29486 49138 29538 49150
rect 16818 49086 16830 49138
rect 16882 49086 16894 49138
rect 22418 49086 22430 49138
rect 22482 49086 22494 49138
rect 26786 49086 26798 49138
rect 26850 49086 26862 49138
rect 11006 49074 11058 49086
rect 20190 49074 20242 49086
rect 24222 49074 24274 49086
rect 29486 49074 29538 49086
rect 30718 49138 30770 49150
rect 30718 49074 30770 49086
rect 32510 49138 32562 49150
rect 32946 49086 32958 49138
rect 33010 49135 33022 49138
rect 33073 49135 33119 49201
rect 33506 49198 33518 49201
rect 33570 49198 33582 49250
rect 38994 49198 39006 49250
rect 39058 49198 39070 49250
rect 33010 49089 33119 49135
rect 36430 49138 36482 49150
rect 33010 49086 33022 49089
rect 32510 49074 32562 49086
rect 36430 49074 36482 49086
rect 37326 49138 37378 49150
rect 37326 49074 37378 49086
rect 39790 49138 39842 49150
rect 39790 49074 39842 49086
rect 41694 49138 41746 49150
rect 41694 49074 41746 49086
rect 43710 49138 43762 49150
rect 43710 49074 43762 49086
rect 44830 49138 44882 49150
rect 44830 49074 44882 49086
rect 53118 49138 53170 49150
rect 53890 49086 53902 49138
rect 53954 49086 53966 49138
rect 57810 49086 57822 49138
rect 57874 49086 57886 49138
rect 53118 49074 53170 49086
rect 7870 49026 7922 49038
rect 9550 49026 9602 49038
rect 4274 48974 4286 49026
rect 4338 48974 4350 49026
rect 7410 48974 7422 49026
rect 7474 48974 7486 49026
rect 9202 48974 9214 49026
rect 9266 48974 9278 49026
rect 7870 48962 7922 48974
rect 9550 48962 9602 48974
rect 9774 49026 9826 49038
rect 13022 49026 13074 49038
rect 19182 49026 19234 49038
rect 24110 49026 24162 49038
rect 27246 49026 27298 49038
rect 11778 48974 11790 49026
rect 11842 48974 11854 49026
rect 12226 48974 12238 49026
rect 12290 48974 12302 49026
rect 12562 48974 12574 49026
rect 12626 48974 12638 49026
rect 13570 48974 13582 49026
rect 13634 48974 13646 49026
rect 13906 48974 13918 49026
rect 13970 48974 13982 49026
rect 14466 48974 14478 49026
rect 14530 48974 14542 49026
rect 15698 48974 15710 49026
rect 15762 48974 15774 49026
rect 16258 48974 16270 49026
rect 16322 48974 16334 49026
rect 16930 48974 16942 49026
rect 16994 48974 17006 49026
rect 17490 48974 17502 49026
rect 17554 48974 17566 49026
rect 19954 48974 19966 49026
rect 20018 48974 20030 49026
rect 21746 48974 21758 49026
rect 21810 48974 21822 49026
rect 22306 48974 22318 49026
rect 22370 48974 22382 49026
rect 23538 48974 23550 49026
rect 23602 48974 23614 49026
rect 26226 48974 26238 49026
rect 26290 48974 26302 49026
rect 9774 48962 9826 48974
rect 13022 48962 13074 48974
rect 19182 48962 19234 48974
rect 24110 48962 24162 48974
rect 27246 48962 27298 48974
rect 28030 49026 28082 49038
rect 28030 48962 28082 48974
rect 28366 49026 28418 49038
rect 28366 48962 28418 48974
rect 28702 49026 28754 49038
rect 29374 49026 29426 49038
rect 29138 48974 29150 49026
rect 29202 48974 29214 49026
rect 28702 48962 28754 48974
rect 29374 48962 29426 48974
rect 33406 49026 33458 49038
rect 33406 48962 33458 48974
rect 37550 49026 37602 49038
rect 37550 48962 37602 48974
rect 38446 49026 38498 49038
rect 38446 48962 38498 48974
rect 39454 49026 39506 49038
rect 39454 48962 39506 48974
rect 39566 49026 39618 49038
rect 39566 48962 39618 48974
rect 40798 49026 40850 49038
rect 43822 49026 43874 49038
rect 41010 48974 41022 49026
rect 41074 48974 41086 49026
rect 40798 48962 40850 48974
rect 43822 48962 43874 48974
rect 46174 49026 46226 49038
rect 46174 48962 46226 48974
rect 47182 49026 47234 49038
rect 47182 48962 47234 48974
rect 53006 49026 53058 49038
rect 53006 48962 53058 48974
rect 53230 49026 53282 49038
rect 54686 49026 54738 49038
rect 54226 48974 54238 49026
rect 54290 48974 54302 49026
rect 55570 48974 55582 49026
rect 55634 48974 55646 49026
rect 53230 48962 53282 48974
rect 54686 48962 54738 48974
rect 8206 48914 8258 48926
rect 8206 48850 8258 48862
rect 10894 48914 10946 48926
rect 27358 48914 27410 48926
rect 14018 48862 14030 48914
rect 14082 48862 14094 48914
rect 17714 48862 17726 48914
rect 17778 48862 17790 48914
rect 22978 48862 22990 48914
rect 23042 48862 23054 48914
rect 10894 48850 10946 48862
rect 27358 48850 27410 48862
rect 29822 48914 29874 48926
rect 29822 48850 29874 48862
rect 31950 48914 32002 48926
rect 38334 48914 38386 48926
rect 37874 48862 37886 48914
rect 37938 48862 37950 48914
rect 31950 48850 32002 48862
rect 38334 48850 38386 48862
rect 38558 48914 38610 48926
rect 38558 48850 38610 48862
rect 39902 48914 39954 48926
rect 39902 48850 39954 48862
rect 43598 48914 43650 48926
rect 43598 48850 43650 48862
rect 44158 48914 44210 48926
rect 44158 48850 44210 48862
rect 45614 48914 45666 48926
rect 45614 48850 45666 48862
rect 45838 48914 45890 48926
rect 45838 48850 45890 48862
rect 46398 48914 46450 48926
rect 46398 48850 46450 48862
rect 46734 48914 46786 48926
rect 46734 48850 46786 48862
rect 51662 48914 51714 48926
rect 51662 48850 51714 48862
rect 51774 48914 51826 48926
rect 51774 48850 51826 48862
rect 4734 48802 4786 48814
rect 4734 48738 4786 48750
rect 11118 48802 11170 48814
rect 11118 48738 11170 48750
rect 15262 48802 15314 48814
rect 15262 48738 15314 48750
rect 27582 48802 27634 48814
rect 27582 48738 27634 48750
rect 27694 48802 27746 48814
rect 27694 48738 27746 48750
rect 27918 48802 27970 48814
rect 27918 48738 27970 48750
rect 28478 48802 28530 48814
rect 28478 48738 28530 48750
rect 29598 48802 29650 48814
rect 29598 48738 29650 48750
rect 30270 48802 30322 48814
rect 30270 48738 30322 48750
rect 31278 48802 31330 48814
rect 31278 48738 31330 48750
rect 31502 48802 31554 48814
rect 31502 48738 31554 48750
rect 31614 48802 31666 48814
rect 31614 48738 31666 48750
rect 31726 48802 31778 48814
rect 31726 48738 31778 48750
rect 32398 48802 32450 48814
rect 32398 48738 32450 48750
rect 32622 48802 32674 48814
rect 32622 48738 32674 48750
rect 32846 48802 32898 48814
rect 32846 48738 32898 48750
rect 34750 48802 34802 48814
rect 34750 48738 34802 48750
rect 40462 48802 40514 48814
rect 40462 48738 40514 48750
rect 44942 48802 44994 48814
rect 44942 48738 44994 48750
rect 45502 48802 45554 48814
rect 45502 48738 45554 48750
rect 47742 48802 47794 48814
rect 47742 48738 47794 48750
rect 51998 48802 52050 48814
rect 51998 48738 52050 48750
rect 52782 48802 52834 48814
rect 52782 48738 52834 48750
rect 1344 48634 58576 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 58576 48634
rect 1344 48548 58576 48582
rect 23326 48466 23378 48478
rect 8082 48414 8094 48466
rect 8146 48414 8158 48466
rect 11554 48414 11566 48466
rect 11618 48414 11630 48466
rect 23326 48402 23378 48414
rect 24222 48466 24274 48478
rect 27470 48466 27522 48478
rect 26786 48414 26798 48466
rect 26850 48414 26862 48466
rect 24222 48402 24274 48414
rect 27470 48402 27522 48414
rect 29374 48466 29426 48478
rect 29374 48402 29426 48414
rect 29822 48466 29874 48478
rect 37102 48466 37154 48478
rect 33058 48414 33070 48466
rect 33122 48414 33134 48466
rect 34514 48414 34526 48466
rect 34578 48414 34590 48466
rect 29822 48402 29874 48414
rect 24670 48354 24722 48366
rect 27582 48354 27634 48366
rect 31502 48354 31554 48366
rect 8978 48302 8990 48354
rect 9042 48302 9054 48354
rect 26114 48302 26126 48354
rect 26178 48302 26190 48354
rect 27682 48302 27694 48354
rect 27746 48302 27758 48354
rect 30594 48302 30606 48354
rect 30658 48302 30670 48354
rect 24670 48290 24722 48302
rect 27582 48290 27634 48302
rect 31502 48290 31554 48302
rect 9886 48242 9938 48254
rect 4274 48190 4286 48242
rect 4338 48190 4350 48242
rect 7970 48190 7982 48242
rect 8034 48190 8046 48242
rect 8754 48190 8766 48242
rect 8818 48190 8830 48242
rect 9886 48178 9938 48190
rect 10446 48242 10498 48254
rect 10446 48178 10498 48190
rect 11230 48242 11282 48254
rect 19294 48242 19346 48254
rect 27246 48242 27298 48254
rect 11330 48190 11342 48242
rect 11394 48190 11406 48242
rect 12450 48190 12462 48242
rect 12514 48190 12526 48242
rect 13458 48190 13470 48242
rect 13522 48190 13534 48242
rect 14802 48190 14814 48242
rect 14866 48190 14878 48242
rect 15250 48190 15262 48242
rect 15314 48190 15326 48242
rect 15586 48190 15598 48242
rect 15650 48190 15662 48242
rect 18610 48190 18622 48242
rect 18674 48190 18686 48242
rect 20066 48190 20078 48242
rect 20130 48190 20142 48242
rect 21074 48190 21086 48242
rect 21138 48190 21150 48242
rect 22306 48190 22318 48242
rect 22370 48190 22382 48242
rect 22866 48190 22878 48242
rect 22930 48190 22942 48242
rect 25778 48190 25790 48242
rect 25842 48190 25854 48242
rect 26786 48190 26798 48242
rect 26850 48190 26862 48242
rect 11230 48178 11282 48190
rect 19294 48178 19346 48190
rect 27246 48178 27298 48190
rect 30270 48242 30322 48254
rect 33073 48242 33119 48414
rect 37102 48402 37154 48414
rect 39006 48466 39058 48478
rect 39006 48402 39058 48414
rect 40126 48466 40178 48478
rect 40126 48402 40178 48414
rect 41022 48466 41074 48478
rect 44270 48466 44322 48478
rect 43474 48414 43486 48466
rect 43538 48414 43550 48466
rect 41022 48402 41074 48414
rect 44270 48402 44322 48414
rect 44830 48466 44882 48478
rect 46162 48414 46174 48466
rect 46226 48414 46238 48466
rect 47058 48414 47070 48466
rect 47122 48414 47134 48466
rect 44830 48402 44882 48414
rect 37998 48354 38050 48366
rect 33618 48302 33630 48354
rect 33682 48302 33694 48354
rect 35074 48302 35086 48354
rect 35138 48302 35150 48354
rect 37762 48302 37774 48354
rect 37826 48302 37838 48354
rect 37998 48290 38050 48302
rect 40910 48354 40962 48366
rect 49422 48354 49474 48366
rect 45154 48302 45166 48354
rect 45218 48302 45230 48354
rect 40910 48290 40962 48302
rect 49422 48290 49474 48302
rect 50878 48354 50930 48366
rect 50878 48290 50930 48302
rect 53230 48354 53282 48366
rect 53230 48290 53282 48302
rect 43822 48242 43874 48254
rect 47406 48242 47458 48254
rect 52446 48242 52498 48254
rect 33058 48190 33070 48242
rect 33122 48190 33134 48242
rect 33506 48190 33518 48242
rect 33570 48190 33582 48242
rect 34402 48190 34414 48242
rect 34466 48190 34478 48242
rect 34962 48190 34974 48242
rect 35026 48190 35038 48242
rect 35970 48190 35982 48242
rect 36034 48190 36046 48242
rect 38210 48190 38222 48242
rect 38274 48190 38286 48242
rect 39890 48190 39902 48242
rect 39954 48190 39966 48242
rect 41234 48190 41246 48242
rect 41298 48190 41310 48242
rect 45490 48190 45502 48242
rect 45554 48190 45566 48242
rect 46050 48190 46062 48242
rect 46114 48190 46126 48242
rect 48962 48190 48974 48242
rect 49026 48190 49038 48242
rect 49186 48190 49198 48242
rect 49250 48190 49262 48242
rect 50306 48190 50318 48242
rect 50370 48190 50382 48242
rect 52098 48190 52110 48242
rect 52162 48190 52174 48242
rect 30270 48178 30322 48190
rect 43822 48178 43874 48190
rect 47406 48178 47458 48190
rect 52446 48178 52498 48190
rect 52670 48242 52722 48254
rect 52670 48178 52722 48190
rect 7646 48130 7698 48142
rect 25454 48130 25506 48142
rect 28366 48130 28418 48142
rect 11554 48078 11566 48130
rect 11618 48078 11630 48130
rect 18498 48078 18510 48130
rect 18562 48078 18574 48130
rect 28018 48078 28030 48130
rect 28082 48078 28094 48130
rect 7646 48066 7698 48078
rect 25454 48066 25506 48078
rect 28366 48066 28418 48078
rect 28590 48130 28642 48142
rect 28590 48066 28642 48078
rect 31054 48130 31106 48142
rect 31054 48066 31106 48078
rect 32062 48130 32114 48142
rect 32062 48066 32114 48078
rect 32622 48130 32674 48142
rect 32622 48066 32674 48078
rect 33182 48130 33234 48142
rect 35758 48130 35810 48142
rect 35522 48078 35534 48130
rect 35586 48078 35598 48130
rect 33182 48066 33234 48078
rect 35758 48066 35810 48078
rect 37662 48130 37714 48142
rect 37662 48066 37714 48078
rect 39454 48130 39506 48142
rect 39454 48066 39506 48078
rect 41694 48130 41746 48142
rect 41694 48066 41746 48078
rect 44158 48130 44210 48142
rect 44158 48066 44210 48078
rect 46734 48130 46786 48142
rect 46734 48066 46786 48078
rect 47742 48130 47794 48142
rect 52558 48130 52610 48142
rect 50082 48078 50094 48130
rect 50146 48078 50158 48130
rect 47742 48066 47794 48078
rect 52558 48066 52610 48078
rect 53118 48130 53170 48142
rect 53118 48066 53170 48078
rect 1934 48018 1986 48030
rect 38670 48018 38722 48030
rect 13458 47966 13470 48018
rect 13522 47966 13534 48018
rect 20626 47966 20638 48018
rect 20690 47966 20702 48018
rect 28914 47966 28926 48018
rect 28978 47966 28990 48018
rect 1934 47954 1986 47966
rect 38670 47954 38722 47966
rect 40238 48018 40290 48030
rect 40238 47954 40290 47966
rect 47854 48018 47906 48030
rect 47854 47954 47906 47966
rect 49534 48018 49586 48030
rect 49534 47954 49586 47966
rect 53006 48018 53058 48030
rect 53006 47954 53058 47966
rect 1344 47850 58576 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 58576 47850
rect 1344 47764 58576 47798
rect 7422 47682 7474 47694
rect 7422 47618 7474 47630
rect 19182 47682 19234 47694
rect 19182 47618 19234 47630
rect 30494 47682 30546 47694
rect 30494 47618 30546 47630
rect 31726 47682 31778 47694
rect 31726 47618 31778 47630
rect 35758 47682 35810 47694
rect 35758 47618 35810 47630
rect 47406 47682 47458 47694
rect 47406 47618 47458 47630
rect 47854 47682 47906 47694
rect 47854 47618 47906 47630
rect 10670 47570 10722 47582
rect 9538 47518 9550 47570
rect 9602 47518 9614 47570
rect 10670 47506 10722 47518
rect 11454 47570 11506 47582
rect 19854 47570 19906 47582
rect 14914 47518 14926 47570
rect 14978 47518 14990 47570
rect 17042 47518 17054 47570
rect 17106 47518 17118 47570
rect 11454 47506 11506 47518
rect 19854 47506 19906 47518
rect 20750 47570 20802 47582
rect 20750 47506 20802 47518
rect 22430 47570 22482 47582
rect 25566 47570 25618 47582
rect 24658 47518 24670 47570
rect 24722 47518 24734 47570
rect 22430 47506 22482 47518
rect 25566 47506 25618 47518
rect 27246 47570 27298 47582
rect 27246 47506 27298 47518
rect 27694 47570 27746 47582
rect 27694 47506 27746 47518
rect 28478 47570 28530 47582
rect 28478 47506 28530 47518
rect 29598 47570 29650 47582
rect 32846 47570 32898 47582
rect 31378 47518 31390 47570
rect 31442 47518 31454 47570
rect 29598 47506 29650 47518
rect 32846 47506 32898 47518
rect 39342 47570 39394 47582
rect 46734 47570 46786 47582
rect 53678 47570 53730 47582
rect 41234 47518 41246 47570
rect 41298 47518 41310 47570
rect 52882 47518 52894 47570
rect 52946 47518 52958 47570
rect 39342 47506 39394 47518
rect 46734 47506 46786 47518
rect 53678 47506 53730 47518
rect 12350 47458 12402 47470
rect 10994 47406 11006 47458
rect 11058 47406 11070 47458
rect 12350 47394 12402 47406
rect 12910 47458 12962 47470
rect 15822 47458 15874 47470
rect 20190 47458 20242 47470
rect 22766 47458 22818 47470
rect 25118 47458 25170 47470
rect 13458 47406 13470 47458
rect 13522 47406 13534 47458
rect 16370 47406 16382 47458
rect 16434 47406 16446 47458
rect 17266 47406 17278 47458
rect 17330 47406 17342 47458
rect 18050 47406 18062 47458
rect 18114 47406 18126 47458
rect 18274 47406 18286 47458
rect 18338 47406 18350 47458
rect 19282 47406 19294 47458
rect 19346 47406 19358 47458
rect 21298 47406 21310 47458
rect 21362 47406 21374 47458
rect 23762 47406 23774 47458
rect 23826 47406 23838 47458
rect 12910 47394 12962 47406
rect 15822 47394 15874 47406
rect 20190 47394 20242 47406
rect 22766 47394 22818 47406
rect 25118 47394 25170 47406
rect 25342 47458 25394 47470
rect 28254 47458 28306 47470
rect 33630 47458 33682 47470
rect 37214 47458 37266 47470
rect 26002 47406 26014 47458
rect 26066 47406 26078 47458
rect 31154 47406 31166 47458
rect 31218 47406 31230 47458
rect 31938 47406 31950 47458
rect 32002 47406 32014 47458
rect 33394 47406 33406 47458
rect 33458 47406 33470 47458
rect 35298 47406 35310 47458
rect 35362 47406 35374 47458
rect 25342 47394 25394 47406
rect 28254 47394 28306 47406
rect 33630 47394 33682 47406
rect 37214 47394 37266 47406
rect 37438 47458 37490 47470
rect 37438 47394 37490 47406
rect 37662 47458 37714 47470
rect 37662 47394 37714 47406
rect 38110 47458 38162 47470
rect 43710 47458 43762 47470
rect 45390 47458 45442 47470
rect 40226 47406 40238 47458
rect 40290 47406 40302 47458
rect 40786 47406 40798 47458
rect 40850 47406 40862 47458
rect 41906 47406 41918 47458
rect 41970 47406 41982 47458
rect 45154 47406 45166 47458
rect 45218 47406 45230 47458
rect 38110 47394 38162 47406
rect 43710 47394 43762 47406
rect 45390 47394 45442 47406
rect 45502 47458 45554 47470
rect 46958 47458 47010 47470
rect 45938 47406 45950 47458
rect 46002 47406 46014 47458
rect 45502 47394 45554 47406
rect 46958 47394 47010 47406
rect 47182 47458 47234 47470
rect 47182 47394 47234 47406
rect 49758 47458 49810 47470
rect 49758 47394 49810 47406
rect 50206 47458 50258 47470
rect 53106 47406 53118 47458
rect 53170 47406 53182 47458
rect 50206 47394 50258 47406
rect 7310 47346 7362 47358
rect 22318 47346 22370 47358
rect 14018 47294 14030 47346
rect 14082 47294 14094 47346
rect 16706 47294 16718 47346
rect 16770 47294 16782 47346
rect 21410 47294 21422 47346
rect 21474 47294 21486 47346
rect 7310 47282 7362 47294
rect 22318 47282 22370 47294
rect 22654 47346 22706 47358
rect 25678 47346 25730 47358
rect 28030 47346 28082 47358
rect 23202 47294 23214 47346
rect 23266 47294 23278 47346
rect 26338 47294 26350 47346
rect 26402 47294 26414 47346
rect 26562 47294 26574 47346
rect 26626 47294 26638 47346
rect 22654 47282 22706 47294
rect 25678 47282 25730 47294
rect 28030 47282 28082 47294
rect 28590 47346 28642 47358
rect 28590 47282 28642 47294
rect 29150 47346 29202 47358
rect 29150 47282 29202 47294
rect 29374 47346 29426 47358
rect 29374 47282 29426 47294
rect 29710 47346 29762 47358
rect 29710 47282 29762 47294
rect 30382 47346 30434 47358
rect 30382 47282 30434 47294
rect 33742 47346 33794 47358
rect 44270 47346 44322 47358
rect 50766 47346 50818 47358
rect 34178 47294 34190 47346
rect 34242 47294 34254 47346
rect 35074 47294 35086 47346
rect 35138 47294 35150 47346
rect 40898 47294 40910 47346
rect 40962 47294 40974 47346
rect 41682 47294 41694 47346
rect 41746 47294 41758 47346
rect 48066 47294 48078 47346
rect 48130 47294 48142 47346
rect 33742 47282 33794 47294
rect 44270 47282 44322 47294
rect 50766 47282 50818 47294
rect 8654 47234 8706 47246
rect 8654 47170 8706 47182
rect 9214 47234 9266 47246
rect 9214 47170 9266 47182
rect 9998 47234 10050 47246
rect 9998 47170 10050 47182
rect 12014 47234 12066 47246
rect 36094 47234 36146 47246
rect 21858 47182 21870 47234
rect 21922 47182 21934 47234
rect 12014 47170 12066 47182
rect 36094 47170 36146 47182
rect 37886 47234 37938 47246
rect 37886 47170 37938 47182
rect 38222 47234 38274 47246
rect 38222 47170 38274 47182
rect 39230 47234 39282 47246
rect 58158 47234 58210 47246
rect 51762 47182 51774 47234
rect 51826 47182 51838 47234
rect 39230 47170 39282 47182
rect 58158 47170 58210 47182
rect 1344 47066 58576 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 58576 47066
rect 1344 46980 58576 47014
rect 11678 46898 11730 46910
rect 11678 46834 11730 46846
rect 13134 46898 13186 46910
rect 13134 46834 13186 46846
rect 13582 46898 13634 46910
rect 13582 46834 13634 46846
rect 16046 46898 16098 46910
rect 18062 46898 18114 46910
rect 16818 46846 16830 46898
rect 16882 46846 16894 46898
rect 16046 46834 16098 46846
rect 18062 46834 18114 46846
rect 20414 46898 20466 46910
rect 20414 46834 20466 46846
rect 20974 46898 21026 46910
rect 20974 46834 21026 46846
rect 29486 46898 29538 46910
rect 29486 46834 29538 46846
rect 33182 46898 33234 46910
rect 33182 46834 33234 46846
rect 35086 46898 35138 46910
rect 35086 46834 35138 46846
rect 38782 46898 38834 46910
rect 40126 46898 40178 46910
rect 39106 46846 39118 46898
rect 39170 46846 39182 46898
rect 38782 46834 38834 46846
rect 40126 46834 40178 46846
rect 40350 46898 40402 46910
rect 50990 46898 51042 46910
rect 45826 46846 45838 46898
rect 45890 46846 45902 46898
rect 53666 46846 53678 46898
rect 53730 46846 53742 46898
rect 40350 46834 40402 46846
rect 50990 46834 51042 46846
rect 6750 46786 6802 46798
rect 6750 46722 6802 46734
rect 8766 46786 8818 46798
rect 11902 46786 11954 46798
rect 9986 46734 9998 46786
rect 10050 46734 10062 46786
rect 10546 46734 10558 46786
rect 10610 46734 10622 46786
rect 11218 46734 11230 46786
rect 11282 46734 11294 46786
rect 8766 46722 8818 46734
rect 11902 46722 11954 46734
rect 14030 46786 14082 46798
rect 14030 46722 14082 46734
rect 14478 46786 14530 46798
rect 14478 46722 14530 46734
rect 14590 46786 14642 46798
rect 14590 46722 14642 46734
rect 16270 46786 16322 46798
rect 16270 46722 16322 46734
rect 21310 46786 21362 46798
rect 21310 46722 21362 46734
rect 27470 46786 27522 46798
rect 27470 46722 27522 46734
rect 29598 46786 29650 46798
rect 29598 46722 29650 46734
rect 29822 46786 29874 46798
rect 34974 46786 35026 46798
rect 30146 46734 30158 46786
rect 30210 46734 30222 46786
rect 29822 46722 29874 46734
rect 34974 46722 35026 46734
rect 35534 46786 35586 46798
rect 39902 46786 39954 46798
rect 45502 46786 45554 46798
rect 36306 46734 36318 46786
rect 36370 46734 36382 46786
rect 41010 46734 41022 46786
rect 41074 46734 41086 46786
rect 44034 46734 44046 46786
rect 44098 46734 44110 46786
rect 35534 46722 35586 46734
rect 39902 46722 39954 46734
rect 45502 46722 45554 46734
rect 48750 46786 48802 46798
rect 48750 46722 48802 46734
rect 49086 46786 49138 46798
rect 49086 46722 49138 46734
rect 50318 46786 50370 46798
rect 52770 46734 52782 46786
rect 52834 46734 52846 46786
rect 50318 46722 50370 46734
rect 7086 46674 7138 46686
rect 12014 46674 12066 46686
rect 9762 46622 9774 46674
rect 9826 46622 9838 46674
rect 10322 46622 10334 46674
rect 10386 46622 10398 46674
rect 7086 46610 7138 46622
rect 12014 46610 12066 46622
rect 12462 46674 12514 46686
rect 12462 46610 12514 46622
rect 17390 46674 17442 46686
rect 18174 46674 18226 46686
rect 17938 46622 17950 46674
rect 18002 46622 18014 46674
rect 17390 46610 17442 46622
rect 18174 46610 18226 46622
rect 18286 46674 18338 46686
rect 18286 46610 18338 46622
rect 18734 46674 18786 46686
rect 19742 46674 19794 46686
rect 18946 46622 18958 46674
rect 19010 46622 19022 46674
rect 18734 46610 18786 46622
rect 19742 46610 19794 46622
rect 20190 46674 20242 46686
rect 20190 46610 20242 46622
rect 22206 46674 22258 46686
rect 28926 46674 28978 46686
rect 22418 46622 22430 46674
rect 22482 46622 22494 46674
rect 22866 46622 22878 46674
rect 22930 46622 22942 46674
rect 23762 46622 23774 46674
rect 23826 46622 23838 46674
rect 27906 46622 27918 46674
rect 27970 46622 27982 46674
rect 22206 46610 22258 46622
rect 28926 46610 28978 46622
rect 29262 46674 29314 46686
rect 35198 46674 35250 46686
rect 40238 46674 40290 46686
rect 44942 46674 44994 46686
rect 30258 46622 30270 46674
rect 30322 46622 30334 46674
rect 32498 46622 32510 46674
rect 32562 46622 32574 46674
rect 35970 46622 35982 46674
rect 36034 46622 36046 46674
rect 36978 46622 36990 46674
rect 37042 46622 37054 46674
rect 40898 46622 40910 46674
rect 40962 46622 40974 46674
rect 41794 46622 41806 46674
rect 41858 46622 41870 46674
rect 42466 46622 42478 46674
rect 42530 46622 42542 46674
rect 42914 46622 42926 46674
rect 42978 46622 42990 46674
rect 29262 46610 29314 46622
rect 35198 46610 35250 46622
rect 40238 46610 40290 46622
rect 44942 46610 44994 46622
rect 45166 46674 45218 46686
rect 48862 46674 48914 46686
rect 46050 46622 46062 46674
rect 46114 46622 46126 46674
rect 45166 46610 45218 46622
rect 48862 46610 48914 46622
rect 49534 46674 49586 46686
rect 49534 46610 49586 46622
rect 50206 46674 50258 46686
rect 51998 46674 52050 46686
rect 50530 46622 50542 46674
rect 50594 46622 50606 46674
rect 51762 46622 51774 46674
rect 51826 46622 51838 46674
rect 50206 46610 50258 46622
rect 51998 46610 52050 46622
rect 52222 46674 52274 46686
rect 52222 46610 52274 46622
rect 52334 46674 52386 46686
rect 52658 46622 52670 46674
rect 52722 46622 52734 46674
rect 53554 46622 53566 46674
rect 53618 46622 53630 46674
rect 52334 46610 52386 46622
rect 11566 46562 11618 46574
rect 11566 46498 11618 46510
rect 16494 46562 16546 46574
rect 16494 46498 16546 46510
rect 20302 46562 20354 46574
rect 20302 46498 20354 46510
rect 21870 46562 21922 46574
rect 25230 46562 25282 46574
rect 24098 46510 24110 46562
rect 24162 46510 24174 46562
rect 21870 46498 21922 46510
rect 25230 46498 25282 46510
rect 26574 46562 26626 46574
rect 26574 46498 26626 46510
rect 27022 46562 27074 46574
rect 27022 46498 27074 46510
rect 28366 46562 28418 46574
rect 34638 46562 34690 46574
rect 31714 46510 31726 46562
rect 31778 46510 31790 46562
rect 28366 46498 28418 46510
rect 34638 46498 34690 46510
rect 36654 46562 36706 46574
rect 36654 46498 36706 46510
rect 36766 46562 36818 46574
rect 36766 46498 36818 46510
rect 37998 46562 38050 46574
rect 37998 46498 38050 46510
rect 38446 46562 38498 46574
rect 45390 46562 45442 46574
rect 41458 46510 41470 46562
rect 41522 46510 41534 46562
rect 38446 46498 38498 46510
rect 45390 46498 45442 46510
rect 49310 46562 49362 46574
rect 49310 46498 49362 46510
rect 49982 46562 50034 46574
rect 49982 46498 50034 46510
rect 8542 46450 8594 46462
rect 8542 46386 8594 46398
rect 8878 46450 8930 46462
rect 8878 46386 8930 46398
rect 14254 46450 14306 46462
rect 14254 46386 14306 46398
rect 14814 46450 14866 46462
rect 14814 46386 14866 46398
rect 15038 46450 15090 46462
rect 15038 46386 15090 46398
rect 17614 46450 17666 46462
rect 21534 46450 21586 46462
rect 25454 46450 25506 46462
rect 19394 46398 19406 46450
rect 19458 46398 19470 46450
rect 20626 46398 20638 46450
rect 20690 46447 20702 46450
rect 21074 46447 21086 46450
rect 20690 46401 21086 46447
rect 20690 46398 20702 46401
rect 21074 46398 21086 46401
rect 21138 46398 21150 46450
rect 23986 46398 23998 46450
rect 24050 46398 24062 46450
rect 25778 46398 25790 46450
rect 25842 46398 25854 46450
rect 17614 46386 17666 46398
rect 21534 46386 21586 46398
rect 25454 46386 25506 46398
rect 1344 46282 58576 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 58576 46282
rect 1344 46196 58576 46230
rect 41246 46114 41298 46126
rect 15698 46062 15710 46114
rect 15762 46062 15774 46114
rect 17602 46062 17614 46114
rect 17666 46062 17678 46114
rect 32834 46062 32846 46114
rect 32898 46062 32910 46114
rect 33842 46062 33854 46114
rect 33906 46111 33918 46114
rect 34626 46111 34638 46114
rect 33906 46065 34638 46111
rect 33906 46062 33918 46065
rect 34626 46062 34638 46065
rect 34690 46062 34702 46114
rect 41246 46050 41298 46062
rect 16382 46002 16434 46014
rect 18734 46002 18786 46014
rect 10322 45950 10334 46002
rect 10386 45950 10398 46002
rect 17490 45950 17502 46002
rect 17554 45950 17566 46002
rect 16382 45938 16434 45950
rect 18734 45938 18786 45950
rect 20302 46002 20354 46014
rect 20302 45938 20354 45950
rect 23102 46002 23154 46014
rect 23102 45938 23154 45950
rect 23886 46002 23938 46014
rect 26238 46002 26290 46014
rect 24770 45950 24782 46002
rect 24834 45950 24846 46002
rect 23886 45938 23938 45950
rect 26238 45938 26290 45950
rect 27358 46002 27410 46014
rect 27358 45938 27410 45950
rect 28590 46002 28642 46014
rect 28590 45938 28642 45950
rect 30046 46002 30098 46014
rect 30046 45938 30098 45950
rect 33854 46002 33906 46014
rect 33854 45938 33906 45950
rect 47966 46002 48018 46014
rect 47966 45938 48018 45950
rect 7198 45890 7250 45902
rect 8094 45890 8146 45902
rect 15598 45890 15650 45902
rect 6066 45838 6078 45890
rect 6130 45838 6142 45890
rect 7634 45838 7646 45890
rect 7698 45838 7710 45890
rect 8866 45838 8878 45890
rect 8930 45838 8942 45890
rect 9538 45838 9550 45890
rect 9602 45838 9614 45890
rect 10098 45838 10110 45890
rect 10162 45838 10174 45890
rect 11778 45838 11790 45890
rect 11842 45838 11854 45890
rect 14130 45838 14142 45890
rect 14194 45838 14206 45890
rect 14354 45838 14366 45890
rect 14418 45838 14430 45890
rect 15474 45838 15486 45890
rect 15538 45838 15550 45890
rect 7198 45826 7250 45838
rect 8094 45826 8146 45838
rect 15598 45826 15650 45838
rect 15934 45890 15986 45902
rect 15934 45826 15986 45838
rect 18958 45890 19010 45902
rect 23774 45890 23826 45902
rect 19170 45838 19182 45890
rect 19234 45838 19246 45890
rect 21298 45838 21310 45890
rect 21362 45838 21374 45890
rect 21858 45838 21870 45890
rect 21922 45838 21934 45890
rect 18958 45826 19010 45838
rect 23774 45826 23826 45838
rect 24670 45890 24722 45902
rect 24670 45826 24722 45838
rect 25678 45890 25730 45902
rect 30158 45890 30210 45902
rect 26562 45838 26574 45890
rect 26626 45838 26638 45890
rect 27682 45838 27694 45890
rect 27746 45838 27758 45890
rect 25678 45826 25730 45838
rect 30158 45826 30210 45838
rect 30382 45890 30434 45902
rect 30382 45826 30434 45838
rect 31278 45890 31330 45902
rect 32286 45890 32338 45902
rect 35422 45890 35474 45902
rect 31490 45838 31502 45890
rect 31554 45838 31566 45890
rect 32386 45838 32398 45890
rect 32450 45838 32462 45890
rect 32722 45838 32734 45890
rect 32786 45838 32798 45890
rect 31278 45826 31330 45838
rect 32286 45826 32338 45838
rect 35422 45826 35474 45838
rect 38558 45890 38610 45902
rect 47406 45890 47458 45902
rect 41570 45838 41582 45890
rect 41634 45838 41646 45890
rect 44930 45838 44942 45890
rect 44994 45838 45006 45890
rect 45266 45838 45278 45890
rect 45330 45838 45342 45890
rect 46050 45838 46062 45890
rect 46114 45838 46126 45890
rect 38558 45826 38610 45838
rect 47406 45826 47458 45838
rect 6302 45778 6354 45790
rect 17838 45778 17890 45790
rect 8754 45726 8766 45778
rect 8818 45726 8830 45778
rect 10434 45726 10446 45778
rect 10498 45726 10510 45778
rect 13458 45726 13470 45778
rect 13522 45726 13534 45778
rect 6302 45714 6354 45726
rect 17838 45714 17890 45726
rect 19742 45778 19794 45790
rect 19742 45714 19794 45726
rect 20190 45778 20242 45790
rect 20190 45714 20242 45726
rect 20526 45778 20578 45790
rect 20526 45714 20578 45726
rect 20750 45778 20802 45790
rect 24110 45778 24162 45790
rect 29150 45778 29202 45790
rect 21970 45726 21982 45778
rect 22034 45726 22046 45778
rect 24434 45726 24446 45778
rect 24498 45726 24510 45778
rect 27010 45726 27022 45778
rect 27074 45726 27086 45778
rect 27346 45726 27358 45778
rect 27410 45726 27422 45778
rect 20750 45714 20802 45726
rect 24110 45714 24162 45726
rect 29150 45714 29202 45726
rect 29262 45778 29314 45790
rect 29262 45714 29314 45726
rect 30494 45778 30546 45790
rect 30494 45714 30546 45726
rect 34862 45778 34914 45790
rect 34862 45714 34914 45726
rect 39006 45778 39058 45790
rect 39006 45714 39058 45726
rect 39230 45778 39282 45790
rect 49646 45778 49698 45790
rect 45490 45726 45502 45778
rect 45554 45726 45566 45778
rect 48738 45726 48750 45778
rect 48802 45726 48814 45778
rect 39230 45714 39282 45726
rect 49646 45714 49698 45726
rect 6638 45666 6690 45678
rect 12910 45666 12962 45678
rect 23438 45666 23490 45678
rect 9426 45614 9438 45666
rect 9490 45614 9502 45666
rect 21522 45614 21534 45666
rect 21586 45614 21598 45666
rect 6638 45602 6690 45614
rect 12910 45602 12962 45614
rect 23438 45602 23490 45614
rect 25118 45666 25170 45678
rect 25118 45602 25170 45614
rect 29486 45666 29538 45678
rect 29486 45602 29538 45614
rect 34302 45666 34354 45678
rect 34302 45602 34354 45614
rect 38782 45666 38834 45678
rect 38782 45602 38834 45614
rect 41358 45666 41410 45678
rect 41358 45602 41410 45614
rect 48414 45666 48466 45678
rect 48414 45602 48466 45614
rect 1344 45498 58576 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 58576 45498
rect 1344 45412 58576 45446
rect 13246 45330 13298 45342
rect 13246 45266 13298 45278
rect 17502 45330 17554 45342
rect 17502 45266 17554 45278
rect 17614 45330 17666 45342
rect 17614 45266 17666 45278
rect 18734 45330 18786 45342
rect 18734 45266 18786 45278
rect 21758 45330 21810 45342
rect 21758 45266 21810 45278
rect 22990 45330 23042 45342
rect 22990 45266 23042 45278
rect 23438 45330 23490 45342
rect 23438 45266 23490 45278
rect 23886 45330 23938 45342
rect 23886 45266 23938 45278
rect 24670 45330 24722 45342
rect 24670 45266 24722 45278
rect 25342 45330 25394 45342
rect 25342 45266 25394 45278
rect 25790 45330 25842 45342
rect 25790 45266 25842 45278
rect 28926 45330 28978 45342
rect 34414 45330 34466 45342
rect 31266 45278 31278 45330
rect 31330 45278 31342 45330
rect 28926 45266 28978 45278
rect 34414 45266 34466 45278
rect 53790 45330 53842 45342
rect 53790 45266 53842 45278
rect 14030 45218 14082 45230
rect 10434 45166 10446 45218
rect 10498 45166 10510 45218
rect 11666 45166 11678 45218
rect 11730 45166 11742 45218
rect 14030 45154 14082 45166
rect 19966 45218 20018 45230
rect 19966 45154 20018 45166
rect 20190 45218 20242 45230
rect 24446 45218 24498 45230
rect 20738 45166 20750 45218
rect 20802 45166 20814 45218
rect 20190 45154 20242 45166
rect 24446 45154 24498 45166
rect 24782 45218 24834 45230
rect 29486 45218 29538 45230
rect 27794 45166 27806 45218
rect 27858 45166 27870 45218
rect 24782 45154 24834 45166
rect 29486 45154 29538 45166
rect 29710 45218 29762 45230
rect 33406 45218 33458 45230
rect 30594 45166 30606 45218
rect 30658 45166 30670 45218
rect 31378 45166 31390 45218
rect 31442 45166 31454 45218
rect 33058 45166 33070 45218
rect 33122 45166 33134 45218
rect 29710 45154 29762 45166
rect 33406 45154 33458 45166
rect 34078 45218 34130 45230
rect 34078 45154 34130 45166
rect 34638 45218 34690 45230
rect 34638 45154 34690 45166
rect 40014 45218 40066 45230
rect 45054 45218 45106 45230
rect 42018 45166 42030 45218
rect 42082 45166 42094 45218
rect 40014 45154 40066 45166
rect 45054 45154 45106 45166
rect 45166 45218 45218 45230
rect 47742 45218 47794 45230
rect 53566 45218 53618 45230
rect 45714 45166 45726 45218
rect 45778 45166 45790 45218
rect 48962 45166 48974 45218
rect 49026 45166 49038 45218
rect 49298 45166 49310 45218
rect 49362 45166 49374 45218
rect 45166 45154 45218 45166
rect 47742 45154 47794 45166
rect 53566 45154 53618 45166
rect 55918 45218 55970 45230
rect 55918 45154 55970 45166
rect 7310 45106 7362 45118
rect 12910 45106 12962 45118
rect 10098 45054 10110 45106
rect 10162 45054 10174 45106
rect 11778 45054 11790 45106
rect 11842 45054 11854 45106
rect 7310 45042 7362 45054
rect 12910 45042 12962 45054
rect 13022 45106 13074 45118
rect 13022 45042 13074 45054
rect 13358 45106 13410 45118
rect 13358 45042 13410 45054
rect 19854 45106 19906 45118
rect 24110 45106 24162 45118
rect 28702 45106 28754 45118
rect 20514 45054 20526 45106
rect 20578 45054 20590 45106
rect 26674 45054 26686 45106
rect 26738 45054 26750 45106
rect 27010 45054 27022 45106
rect 27074 45054 27086 45106
rect 27906 45054 27918 45106
rect 27970 45054 27982 45106
rect 28466 45054 28478 45106
rect 28530 45054 28542 45106
rect 19854 45042 19906 45054
rect 24110 45042 24162 45054
rect 28702 45042 28754 45054
rect 28814 45106 28866 45118
rect 34302 45106 34354 45118
rect 45278 45106 45330 45118
rect 29138 45054 29150 45106
rect 29202 45054 29214 45106
rect 30706 45054 30718 45106
rect 30770 45054 30782 45106
rect 31154 45054 31166 45106
rect 31218 45054 31230 45106
rect 32498 45054 32510 45106
rect 32562 45054 32574 45106
rect 35298 45054 35310 45106
rect 35362 45054 35374 45106
rect 35522 45054 35534 45106
rect 35586 45054 35598 45106
rect 36194 45054 36206 45106
rect 36258 45054 36270 45106
rect 40338 45054 40350 45106
rect 40402 45054 40414 45106
rect 41346 45054 41358 45106
rect 41410 45054 41422 45106
rect 42130 45054 42142 45106
rect 42194 45054 42206 45106
rect 28814 45042 28866 45054
rect 34302 45042 34354 45054
rect 45278 45042 45330 45054
rect 46846 45106 46898 45118
rect 46846 45042 46898 45054
rect 47070 45106 47122 45118
rect 55246 45106 55298 45118
rect 48738 45054 48750 45106
rect 48802 45054 48814 45106
rect 50306 45054 50318 45106
rect 50370 45054 50382 45106
rect 50978 45054 50990 45106
rect 51042 45054 51054 45106
rect 54562 45054 54574 45106
rect 54626 45054 54638 45106
rect 47070 45042 47122 45054
rect 55246 45042 55298 45054
rect 55582 45106 55634 45118
rect 55582 45042 55634 45054
rect 7870 44994 7922 45006
rect 14926 44994 14978 45006
rect 14130 44942 14142 44994
rect 14194 44942 14206 44994
rect 7870 44930 7922 44942
rect 14926 44930 14978 44942
rect 15262 44994 15314 45006
rect 15262 44930 15314 44942
rect 15710 44994 15762 45006
rect 15710 44930 15762 44942
rect 16382 44994 16434 45006
rect 16382 44930 16434 44942
rect 16830 44994 16882 45006
rect 16830 44930 16882 44942
rect 18286 44994 18338 45006
rect 18286 44930 18338 44942
rect 19070 44994 19122 45006
rect 19070 44930 19122 44942
rect 19518 44994 19570 45006
rect 19518 44930 19570 44942
rect 21198 44994 21250 45006
rect 21198 44930 21250 44942
rect 22094 44994 22146 45006
rect 22094 44930 22146 44942
rect 26238 44994 26290 45006
rect 29598 44994 29650 45006
rect 28018 44942 28030 44994
rect 28082 44942 28094 44994
rect 26238 44930 26290 44942
rect 29598 44930 29650 44942
rect 38334 44994 38386 45006
rect 46622 44994 46674 45006
rect 41794 44942 41806 44994
rect 41858 44942 41870 44994
rect 38334 44930 38386 44942
rect 46622 44930 46674 44942
rect 49982 44994 50034 45006
rect 50754 44942 50766 44994
rect 50818 44942 50830 44994
rect 53890 44942 53902 44994
rect 53954 44942 53966 44994
rect 54338 44942 54350 44994
rect 54402 44942 54414 44994
rect 49982 44930 50034 44942
rect 13806 44882 13858 44894
rect 13806 44818 13858 44830
rect 17726 44882 17778 44894
rect 17726 44818 17778 44830
rect 36430 44882 36482 44894
rect 36430 44818 36482 44830
rect 40350 44882 40402 44894
rect 40350 44818 40402 44830
rect 47294 44882 47346 44894
rect 51202 44830 51214 44882
rect 51266 44830 51278 44882
rect 47294 44818 47346 44830
rect 1344 44714 58576 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 58576 44714
rect 1344 44628 58576 44662
rect 7534 44546 7586 44558
rect 7534 44482 7586 44494
rect 14814 44546 14866 44558
rect 14814 44482 14866 44494
rect 19294 44546 19346 44558
rect 29262 44546 29314 44558
rect 24882 44494 24894 44546
rect 24946 44494 24958 44546
rect 19294 44482 19346 44494
rect 29262 44482 29314 44494
rect 30046 44546 30098 44558
rect 30046 44482 30098 44494
rect 43374 44546 43426 44558
rect 43374 44482 43426 44494
rect 43486 44546 43538 44558
rect 43486 44482 43538 44494
rect 46734 44546 46786 44558
rect 46734 44482 46786 44494
rect 46958 44546 47010 44558
rect 46958 44482 47010 44494
rect 47406 44546 47458 44558
rect 47406 44482 47458 44494
rect 47518 44546 47570 44558
rect 47518 44482 47570 44494
rect 22318 44434 22370 44446
rect 16706 44382 16718 44434
rect 16770 44382 16782 44434
rect 16930 44382 16942 44434
rect 16994 44382 17006 44434
rect 18834 44382 18846 44434
rect 18898 44382 18910 44434
rect 22318 44370 22370 44382
rect 23998 44434 24050 44446
rect 23998 44370 24050 44382
rect 28590 44434 28642 44446
rect 34526 44434 34578 44446
rect 38222 44434 38274 44446
rect 32610 44382 32622 44434
rect 32674 44382 32686 44434
rect 37874 44382 37886 44434
rect 37938 44382 37950 44434
rect 28590 44370 28642 44382
rect 34526 44370 34578 44382
rect 38222 44370 38274 44382
rect 39230 44434 39282 44446
rect 39230 44370 39282 44382
rect 39342 44434 39394 44446
rect 49310 44434 49362 44446
rect 51326 44434 51378 44446
rect 57934 44434 57986 44446
rect 41346 44382 41358 44434
rect 41410 44382 41422 44434
rect 50866 44382 50878 44434
rect 50930 44382 50942 44434
rect 53666 44382 53678 44434
rect 53730 44382 53742 44434
rect 54674 44382 54686 44434
rect 54738 44382 54750 44434
rect 39342 44370 39394 44382
rect 49310 44370 49362 44382
rect 51326 44370 51378 44382
rect 57934 44370 57986 44382
rect 9998 44322 10050 44334
rect 9998 44258 10050 44270
rect 12910 44322 12962 44334
rect 12910 44258 12962 44270
rect 15710 44322 15762 44334
rect 19854 44322 19906 44334
rect 16594 44270 16606 44322
rect 16658 44270 16670 44322
rect 17266 44270 17278 44322
rect 17330 44270 17342 44322
rect 18498 44270 18510 44322
rect 18562 44270 18574 44322
rect 19058 44270 19070 44322
rect 19122 44270 19134 44322
rect 15710 44258 15762 44270
rect 19854 44258 19906 44270
rect 21310 44322 21362 44334
rect 21310 44258 21362 44270
rect 21870 44322 21922 44334
rect 21870 44258 21922 44270
rect 23886 44322 23938 44334
rect 23886 44258 23938 44270
rect 24110 44322 24162 44334
rect 24110 44258 24162 44270
rect 24558 44322 24610 44334
rect 26462 44322 26514 44334
rect 29486 44322 29538 44334
rect 24994 44270 25006 44322
rect 25058 44270 25070 44322
rect 26786 44270 26798 44322
rect 26850 44270 26862 44322
rect 24558 44258 24610 44270
rect 26462 44258 26514 44270
rect 29486 44258 29538 44270
rect 29710 44322 29762 44334
rect 29710 44258 29762 44270
rect 30606 44322 30658 44334
rect 35982 44322 36034 44334
rect 41022 44322 41074 44334
rect 31826 44270 31838 44322
rect 31890 44270 31902 44322
rect 32274 44270 32286 44322
rect 32338 44270 32350 44322
rect 32834 44270 32846 44322
rect 32898 44270 32910 44322
rect 33954 44270 33966 44322
rect 34018 44270 34030 44322
rect 34962 44270 34974 44322
rect 35026 44270 35038 44322
rect 37538 44270 37550 44322
rect 37602 44270 37614 44322
rect 38994 44270 39006 44322
rect 39058 44270 39070 44322
rect 39666 44270 39678 44322
rect 39730 44270 39742 44322
rect 40786 44270 40798 44322
rect 40850 44270 40862 44322
rect 30606 44258 30658 44270
rect 35982 44258 36034 44270
rect 41022 44258 41074 44270
rect 41246 44322 41298 44334
rect 42702 44322 42754 44334
rect 41458 44270 41470 44322
rect 41522 44270 41534 44322
rect 41246 44258 41298 44270
rect 42702 44258 42754 44270
rect 43150 44322 43202 44334
rect 43150 44258 43202 44270
rect 45054 44322 45106 44334
rect 47294 44322 47346 44334
rect 45378 44270 45390 44322
rect 45442 44270 45454 44322
rect 45826 44270 45838 44322
rect 45890 44270 45902 44322
rect 48850 44270 48862 44322
rect 48914 44270 48926 44322
rect 50642 44270 50654 44322
rect 50706 44270 50718 44322
rect 53778 44270 53790 44322
rect 53842 44270 53854 44322
rect 54562 44270 54574 44322
rect 54626 44270 54638 44322
rect 55906 44270 55918 44322
rect 55970 44270 55982 44322
rect 45054 44258 45106 44270
rect 47294 44258 47346 44270
rect 7310 44210 7362 44222
rect 7310 44146 7362 44158
rect 14478 44210 14530 44222
rect 19966 44210 20018 44222
rect 17602 44158 17614 44210
rect 17666 44158 17678 44210
rect 14478 44146 14530 44158
rect 19966 44146 20018 44158
rect 20526 44210 20578 44222
rect 29822 44210 29874 44222
rect 25330 44158 25342 44210
rect 25394 44158 25406 44210
rect 20526 44146 20578 44158
rect 29822 44146 29874 44158
rect 31054 44210 31106 44222
rect 31054 44146 31106 44158
rect 31278 44210 31330 44222
rect 35646 44210 35698 44222
rect 33058 44158 33070 44210
rect 33122 44158 33134 44210
rect 33842 44158 33854 44210
rect 33906 44158 33918 44210
rect 34514 44158 34526 44210
rect 34578 44158 34590 44210
rect 38770 44158 38782 44210
rect 38834 44158 38846 44210
rect 54898 44158 54910 44210
rect 54962 44158 54974 44210
rect 31278 44146 31330 44158
rect 35646 44146 35698 44158
rect 7870 44098 7922 44110
rect 7870 44034 7922 44046
rect 10110 44098 10162 44110
rect 10110 44034 10162 44046
rect 10334 44098 10386 44110
rect 10334 44034 10386 44046
rect 12350 44098 12402 44110
rect 12350 44034 12402 44046
rect 13582 44098 13634 44110
rect 13582 44034 13634 44046
rect 14030 44098 14082 44110
rect 14030 44034 14082 44046
rect 14702 44098 14754 44110
rect 14702 44034 14754 44046
rect 15150 44098 15202 44110
rect 15150 44034 15202 44046
rect 20190 44098 20242 44110
rect 20190 44034 20242 44046
rect 23102 44098 23154 44110
rect 23102 44034 23154 44046
rect 23550 44098 23602 44110
rect 23550 44034 23602 44046
rect 30942 44098 30994 44110
rect 30942 44034 30994 44046
rect 35758 44098 35810 44110
rect 35758 44034 35810 44046
rect 36318 44098 36370 44110
rect 36318 44034 36370 44046
rect 43486 44098 43538 44110
rect 43486 44034 43538 44046
rect 44830 44098 44882 44110
rect 44830 44034 44882 44046
rect 44942 44098 44994 44110
rect 46050 44046 46062 44098
rect 46114 44046 46126 44098
rect 44942 44034 44994 44046
rect 1344 43930 58576 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 58576 43930
rect 1344 43844 58576 43878
rect 29934 43762 29986 43774
rect 6962 43710 6974 43762
rect 7026 43710 7038 43762
rect 8082 43710 8094 43762
rect 8146 43710 8158 43762
rect 29934 43698 29986 43710
rect 33406 43762 33458 43774
rect 33406 43698 33458 43710
rect 33742 43762 33794 43774
rect 33742 43698 33794 43710
rect 34414 43762 34466 43774
rect 34414 43698 34466 43710
rect 41246 43762 41298 43774
rect 41246 43698 41298 43710
rect 46734 43762 46786 43774
rect 46734 43698 46786 43710
rect 49870 43762 49922 43774
rect 49870 43698 49922 43710
rect 54126 43762 54178 43774
rect 54126 43698 54178 43710
rect 7646 43650 7698 43662
rect 14926 43650 14978 43662
rect 23214 43650 23266 43662
rect 14354 43598 14366 43650
rect 14418 43598 14430 43650
rect 18386 43598 18398 43650
rect 18450 43598 18462 43650
rect 21074 43598 21086 43650
rect 21138 43598 21150 43650
rect 7646 43586 7698 43598
rect 14926 43586 14978 43598
rect 23214 43586 23266 43598
rect 23438 43650 23490 43662
rect 23438 43586 23490 43598
rect 24334 43650 24386 43662
rect 24334 43586 24386 43598
rect 27022 43650 27074 43662
rect 27022 43586 27074 43598
rect 29038 43650 29090 43662
rect 29038 43586 29090 43598
rect 29150 43650 29202 43662
rect 29150 43586 29202 43598
rect 30830 43650 30882 43662
rect 30830 43586 30882 43598
rect 31390 43650 31442 43662
rect 31390 43586 31442 43598
rect 34638 43650 34690 43662
rect 34638 43586 34690 43598
rect 36654 43650 36706 43662
rect 36654 43586 36706 43598
rect 36766 43650 36818 43662
rect 36766 43586 36818 43598
rect 51438 43650 51490 43662
rect 51438 43586 51490 43598
rect 53118 43650 53170 43662
rect 53118 43586 53170 43598
rect 53902 43650 53954 43662
rect 53902 43586 53954 43598
rect 56590 43650 56642 43662
rect 56590 43586 56642 43598
rect 6638 43538 6690 43550
rect 6638 43474 6690 43486
rect 7422 43538 7474 43550
rect 7422 43474 7474 43486
rect 7534 43538 7586 43550
rect 14814 43538 14866 43550
rect 23774 43538 23826 43550
rect 28030 43538 28082 43550
rect 9538 43486 9550 43538
rect 9602 43486 9614 43538
rect 11106 43486 11118 43538
rect 11170 43486 11182 43538
rect 12338 43486 12350 43538
rect 12402 43486 12414 43538
rect 13346 43486 13358 43538
rect 13410 43486 13422 43538
rect 13906 43486 13918 43538
rect 13970 43486 13982 43538
rect 16146 43486 16158 43538
rect 16210 43486 16222 43538
rect 17714 43486 17726 43538
rect 17778 43486 17790 43538
rect 18162 43486 18174 43538
rect 18226 43486 18238 43538
rect 18946 43486 18958 43538
rect 19010 43486 19022 43538
rect 19506 43486 19518 43538
rect 19570 43486 19582 43538
rect 20402 43486 20414 43538
rect 20466 43486 20478 43538
rect 20962 43486 20974 43538
rect 21026 43486 21038 43538
rect 21858 43486 21870 43538
rect 21922 43486 21934 43538
rect 25330 43486 25342 43538
rect 25394 43486 25406 43538
rect 25554 43486 25566 43538
rect 25618 43486 25630 43538
rect 26562 43486 26574 43538
rect 26626 43486 26638 43538
rect 7534 43474 7586 43486
rect 14814 43474 14866 43486
rect 23774 43474 23826 43486
rect 28030 43474 28082 43486
rect 29598 43538 29650 43550
rect 29598 43474 29650 43486
rect 30382 43538 30434 43550
rect 30382 43474 30434 43486
rect 34862 43538 34914 43550
rect 40910 43538 40962 43550
rect 44382 43538 44434 43550
rect 51326 43538 51378 43550
rect 36418 43486 36430 43538
rect 36482 43486 36494 43538
rect 37762 43486 37774 43538
rect 37826 43486 37838 43538
rect 42578 43486 42590 43538
rect 42642 43486 42654 43538
rect 43698 43486 43710 43538
rect 43762 43486 43774 43538
rect 45266 43486 45278 43538
rect 45330 43486 45342 43538
rect 49074 43486 49086 43538
rect 49138 43486 49150 43538
rect 34862 43474 34914 43486
rect 40910 43474 40962 43486
rect 44382 43474 44434 43486
rect 51326 43474 51378 43486
rect 51662 43538 51714 43550
rect 53454 43538 53506 43550
rect 55470 43538 55522 43550
rect 52210 43486 52222 43538
rect 52274 43486 52286 43538
rect 54786 43486 54798 43538
rect 54850 43486 54862 43538
rect 56802 43486 56814 43538
rect 56866 43486 56878 43538
rect 51662 43474 51714 43486
rect 53454 43474 53506 43486
rect 55470 43474 55522 43486
rect 15710 43426 15762 43438
rect 17390 43426 17442 43438
rect 22766 43426 22818 43438
rect 10322 43374 10334 43426
rect 10386 43374 10398 43426
rect 16482 43374 16494 43426
rect 16546 43374 16558 43426
rect 21634 43374 21646 43426
rect 21698 43374 21710 43426
rect 15710 43362 15762 43374
rect 17390 43362 17442 43374
rect 22766 43362 22818 43374
rect 27694 43426 27746 43438
rect 27694 43362 27746 43374
rect 34750 43426 34802 43438
rect 38558 43426 38610 43438
rect 38434 43374 38446 43426
rect 38498 43374 38510 43426
rect 34750 43362 34802 43374
rect 38558 43362 38610 43374
rect 46174 43426 46226 43438
rect 46174 43362 46226 43374
rect 49310 43426 49362 43438
rect 54014 43426 54066 43438
rect 52322 43374 52334 43426
rect 52386 43374 52398 43426
rect 54562 43374 54574 43426
rect 54626 43374 54638 43426
rect 49310 43362 49362 43374
rect 54014 43362 54066 43374
rect 11118 43314 11170 43326
rect 11118 43250 11170 43262
rect 11454 43314 11506 43326
rect 11454 43250 11506 43262
rect 14926 43314 14978 43326
rect 14926 43250 14978 43262
rect 23102 43314 23154 43326
rect 23102 43250 23154 43262
rect 26462 43314 26514 43326
rect 26462 43250 26514 43262
rect 28254 43314 28306 43326
rect 29038 43314 29090 43326
rect 49422 43314 49474 43326
rect 28578 43262 28590 43314
rect 28642 43262 28654 43314
rect 37202 43262 37214 43314
rect 37266 43262 37278 43314
rect 45266 43262 45278 43314
rect 45330 43262 45342 43314
rect 28254 43250 28306 43262
rect 29038 43250 29090 43262
rect 49422 43250 49474 43262
rect 1344 43146 58576 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 58576 43146
rect 1344 43060 58576 43094
rect 29598 42978 29650 42990
rect 16594 42926 16606 42978
rect 16658 42926 16670 42978
rect 18722 42926 18734 42978
rect 18786 42926 18798 42978
rect 28018 42926 28030 42978
rect 28082 42926 28094 42978
rect 29598 42914 29650 42926
rect 30718 42978 30770 42990
rect 57934 42978 57986 42990
rect 36306 42926 36318 42978
rect 36370 42926 36382 42978
rect 45826 42926 45838 42978
rect 45890 42926 45902 42978
rect 30718 42914 30770 42926
rect 57934 42914 57986 42926
rect 1710 42866 1762 42878
rect 12126 42866 12178 42878
rect 7634 42814 7646 42866
rect 7698 42814 7710 42866
rect 1710 42802 1762 42814
rect 12126 42802 12178 42814
rect 12686 42866 12738 42878
rect 21534 42866 21586 42878
rect 29822 42866 29874 42878
rect 37774 42866 37826 42878
rect 51214 42866 51266 42878
rect 53678 42866 53730 42878
rect 18274 42814 18286 42866
rect 18338 42814 18350 42866
rect 19506 42814 19518 42866
rect 19570 42814 19582 42866
rect 26562 42814 26574 42866
rect 26626 42814 26638 42866
rect 27458 42814 27470 42866
rect 27522 42814 27534 42866
rect 34402 42814 34414 42866
rect 34466 42814 34478 42866
rect 38434 42814 38446 42866
rect 38498 42814 38510 42866
rect 42914 42814 42926 42866
rect 42978 42814 42990 42866
rect 45378 42814 45390 42866
rect 45442 42814 45454 42866
rect 52770 42814 52782 42866
rect 52834 42814 52846 42866
rect 12686 42802 12738 42814
rect 21534 42802 21586 42814
rect 29822 42802 29874 42814
rect 37774 42802 37826 42814
rect 51214 42802 51266 42814
rect 53678 42802 53730 42814
rect 21310 42754 21362 42766
rect 7298 42702 7310 42754
rect 7362 42702 7374 42754
rect 7858 42702 7870 42754
rect 7922 42702 7934 42754
rect 10322 42702 10334 42754
rect 10386 42702 10398 42754
rect 13794 42702 13806 42754
rect 13858 42702 13870 42754
rect 15026 42702 15038 42754
rect 15090 42702 15102 42754
rect 16034 42702 16046 42754
rect 16098 42702 16110 42754
rect 17602 42702 17614 42754
rect 17666 42702 17678 42754
rect 18722 42702 18734 42754
rect 18786 42702 18798 42754
rect 19730 42702 19742 42754
rect 19794 42702 19806 42754
rect 20514 42702 20526 42754
rect 20578 42702 20590 42754
rect 21310 42690 21362 42702
rect 22318 42754 22370 42766
rect 28702 42754 28754 42766
rect 22978 42702 22990 42754
rect 23042 42702 23054 42754
rect 24434 42702 24446 42754
rect 24498 42702 24510 42754
rect 25890 42702 25902 42754
rect 25954 42702 25966 42754
rect 26786 42702 26798 42754
rect 26850 42702 26862 42754
rect 27570 42702 27582 42754
rect 27634 42702 27646 42754
rect 22318 42690 22370 42702
rect 28702 42690 28754 42702
rect 29038 42754 29090 42766
rect 29038 42690 29090 42702
rect 30382 42754 30434 42766
rect 30382 42690 30434 42702
rect 31838 42754 31890 42766
rect 31838 42690 31890 42702
rect 32398 42754 32450 42766
rect 37438 42754 37490 42766
rect 34290 42702 34302 42754
rect 34354 42702 34366 42754
rect 36082 42702 36094 42754
rect 36146 42702 36158 42754
rect 32398 42690 32450 42702
rect 37438 42690 37490 42702
rect 37550 42754 37602 42766
rect 41358 42754 41410 42766
rect 38546 42702 38558 42754
rect 38610 42702 38622 42754
rect 37550 42690 37602 42702
rect 41358 42690 41410 42702
rect 41918 42754 41970 42766
rect 47966 42754 48018 42766
rect 42242 42702 42254 42754
rect 42306 42702 42318 42754
rect 44930 42702 44942 42754
rect 44994 42702 45006 42754
rect 45490 42702 45502 42754
rect 45554 42702 45566 42754
rect 41918 42690 41970 42702
rect 47966 42690 48018 42702
rect 48190 42754 48242 42766
rect 48190 42690 48242 42702
rect 48414 42754 48466 42766
rect 49410 42702 49422 42754
rect 49474 42702 49486 42754
rect 52994 42702 53006 42754
rect 53058 42702 53070 42754
rect 56018 42702 56030 42754
rect 56082 42702 56094 42754
rect 48414 42690 48466 42702
rect 9774 42642 9826 42654
rect 8306 42590 8318 42642
rect 8370 42590 8382 42642
rect 9774 42578 9826 42590
rect 10894 42642 10946 42654
rect 30046 42642 30098 42654
rect 16258 42590 16270 42642
rect 16322 42590 16334 42642
rect 19394 42590 19406 42642
rect 19458 42590 19470 42642
rect 24882 42590 24894 42642
rect 24946 42590 24958 42642
rect 26002 42590 26014 42642
rect 26066 42590 26078 42642
rect 29362 42590 29374 42642
rect 29426 42590 29438 42642
rect 10894 42578 10946 42590
rect 30046 42578 30098 42590
rect 31502 42642 31554 42654
rect 31502 42578 31554 42590
rect 32510 42642 32562 42654
rect 32510 42578 32562 42590
rect 32734 42642 32786 42654
rect 37886 42642 37938 42654
rect 35522 42590 35534 42642
rect 35586 42590 35598 42642
rect 32734 42578 32786 42590
rect 37886 42578 37938 42590
rect 38222 42642 38274 42654
rect 49982 42642 50034 42654
rect 42578 42590 42590 42642
rect 42642 42590 42654 42642
rect 38222 42578 38274 42590
rect 49982 42578 50034 42590
rect 9214 42530 9266 42542
rect 30158 42530 30210 42542
rect 21858 42478 21870 42530
rect 21922 42478 21934 42530
rect 24098 42478 24110 42530
rect 24162 42478 24174 42530
rect 9214 42466 9266 42478
rect 30158 42466 30210 42478
rect 30606 42530 30658 42542
rect 30606 42466 30658 42478
rect 31166 42530 31218 42542
rect 31166 42466 31218 42478
rect 31614 42530 31666 42542
rect 31614 42466 31666 42478
rect 39006 42530 39058 42542
rect 39006 42466 39058 42478
rect 48862 42530 48914 42542
rect 48862 42466 48914 42478
rect 50878 42530 50930 42542
rect 50878 42466 50930 42478
rect 1344 42362 58576 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 58576 42362
rect 1344 42276 58576 42310
rect 21646 42194 21698 42206
rect 30270 42194 30322 42206
rect 8530 42142 8542 42194
rect 8594 42142 8606 42194
rect 13906 42142 13918 42194
rect 13970 42142 13982 42194
rect 27906 42142 27918 42194
rect 27970 42142 27982 42194
rect 21646 42130 21698 42142
rect 30270 42130 30322 42142
rect 30830 42194 30882 42206
rect 30830 42130 30882 42142
rect 33182 42194 33234 42206
rect 33182 42130 33234 42142
rect 33742 42194 33794 42206
rect 33742 42130 33794 42142
rect 41358 42194 41410 42206
rect 41358 42130 41410 42142
rect 42366 42194 42418 42206
rect 42366 42130 42418 42142
rect 46510 42194 46562 42206
rect 46510 42130 46562 42142
rect 49086 42194 49138 42206
rect 49086 42130 49138 42142
rect 51550 42194 51602 42206
rect 51550 42130 51602 42142
rect 51774 42194 51826 42206
rect 51774 42130 51826 42142
rect 52558 42194 52610 42206
rect 52558 42130 52610 42142
rect 10782 42082 10834 42094
rect 10782 42018 10834 42030
rect 12574 42082 12626 42094
rect 12574 42018 12626 42030
rect 13470 42082 13522 42094
rect 13470 42018 13522 42030
rect 15486 42082 15538 42094
rect 15486 42018 15538 42030
rect 19630 42082 19682 42094
rect 23662 42082 23714 42094
rect 19954 42030 19966 42082
rect 20018 42030 20030 42082
rect 20738 42030 20750 42082
rect 20802 42030 20814 42082
rect 22978 42030 22990 42082
rect 23042 42030 23054 42082
rect 19630 42018 19682 42030
rect 23662 42018 23714 42030
rect 25566 42082 25618 42094
rect 28926 42082 28978 42094
rect 27458 42030 27470 42082
rect 27522 42030 27534 42082
rect 28130 42030 28142 42082
rect 28194 42030 28206 42082
rect 25566 42018 25618 42030
rect 28926 42018 28978 42030
rect 29150 42082 29202 42094
rect 29150 42018 29202 42030
rect 31054 42082 31106 42094
rect 31054 42018 31106 42030
rect 34862 42082 34914 42094
rect 34862 42018 34914 42030
rect 35086 42082 35138 42094
rect 35086 42018 35138 42030
rect 35646 42082 35698 42094
rect 35646 42018 35698 42030
rect 47518 42082 47570 42094
rect 47518 42018 47570 42030
rect 49310 42082 49362 42094
rect 49310 42018 49362 42030
rect 11342 41970 11394 41982
rect 14590 41970 14642 41982
rect 19406 41970 19458 41982
rect 12114 41918 12126 41970
rect 12178 41918 12190 41970
rect 12450 41918 12462 41970
rect 12514 41918 12526 41970
rect 14914 41918 14926 41970
rect 14978 41918 14990 41970
rect 17378 41918 17390 41970
rect 17442 41918 17454 41970
rect 18274 41918 18286 41970
rect 18338 41918 18350 41970
rect 11342 41906 11394 41918
rect 14590 41906 14642 41918
rect 19406 41906 19458 41918
rect 19742 41970 19794 41982
rect 19742 41906 19794 41918
rect 21422 41970 21474 41982
rect 21422 41906 21474 41918
rect 21534 41970 21586 41982
rect 21534 41906 21586 41918
rect 21870 41970 21922 41982
rect 21870 41906 21922 41918
rect 22654 41970 22706 41982
rect 25342 41970 25394 41982
rect 29822 41970 29874 41982
rect 22866 41918 22878 41970
rect 22930 41918 22942 41970
rect 23874 41918 23886 41970
rect 23938 41918 23950 41970
rect 26450 41918 26462 41970
rect 26514 41918 26526 41970
rect 27346 41918 27358 41970
rect 27410 41918 27422 41970
rect 28466 41918 28478 41970
rect 28530 41918 28542 41970
rect 29362 41918 29374 41970
rect 29426 41918 29438 41970
rect 22654 41906 22706 41918
rect 25342 41906 25394 41918
rect 29822 41906 29874 41918
rect 30494 41970 30546 41982
rect 30494 41906 30546 41918
rect 31166 41970 31218 41982
rect 31166 41906 31218 41918
rect 34190 41970 34242 41982
rect 35198 41970 35250 41982
rect 39790 41970 39842 41982
rect 34626 41918 34638 41970
rect 34690 41918 34702 41970
rect 35858 41918 35870 41970
rect 35922 41918 35934 41970
rect 34190 41906 34242 41918
rect 35198 41906 35250 41918
rect 39790 41906 39842 41918
rect 42142 41970 42194 41982
rect 42142 41906 42194 41918
rect 42478 41970 42530 41982
rect 45726 41970 45778 41982
rect 45266 41918 45278 41970
rect 45330 41918 45342 41970
rect 42478 41906 42530 41918
rect 45726 41906 45778 41918
rect 45950 41970 46002 41982
rect 47294 41970 47346 41982
rect 46274 41918 46286 41970
rect 46338 41918 46350 41970
rect 45950 41906 46002 41918
rect 47294 41906 47346 41918
rect 47742 41970 47794 41982
rect 47742 41906 47794 41918
rect 47854 41970 47906 41982
rect 49198 41970 49250 41982
rect 48738 41918 48750 41970
rect 48802 41918 48814 41970
rect 47854 41906 47906 41918
rect 49198 41906 49250 41918
rect 49758 41970 49810 41982
rect 51214 41970 51266 41982
rect 50082 41918 50094 41970
rect 50146 41918 50158 41970
rect 49758 41906 49810 41918
rect 51214 41906 51266 41918
rect 51886 41970 51938 41982
rect 51886 41906 51938 41918
rect 52446 41970 52498 41982
rect 52446 41906 52498 41918
rect 52782 41970 52834 41982
rect 52782 41906 52834 41918
rect 7982 41858 8034 41870
rect 22094 41858 22146 41870
rect 29262 41858 29314 41870
rect 17938 41806 17950 41858
rect 18002 41806 18014 41858
rect 25666 41806 25678 41858
rect 25730 41806 25742 41858
rect 7982 41794 8034 41806
rect 22094 41794 22146 41806
rect 29262 41794 29314 41806
rect 34974 41858 35026 41870
rect 41918 41858 41970 41870
rect 40226 41806 40238 41858
rect 40290 41806 40302 41858
rect 34974 41794 35026 41806
rect 41918 41794 41970 41806
rect 44382 41858 44434 41870
rect 50654 41858 50706 41870
rect 44818 41806 44830 41858
rect 44882 41806 44894 41858
rect 44382 41794 44434 41806
rect 50654 41794 50706 41806
rect 8206 41746 8258 41758
rect 22318 41746 22370 41758
rect 46174 41746 46226 41758
rect 18386 41694 18398 41746
rect 18450 41694 18462 41746
rect 29586 41694 29598 41746
rect 29650 41743 29662 41746
rect 30258 41743 30270 41746
rect 29650 41697 30270 41743
rect 29650 41694 29662 41697
rect 30258 41694 30270 41697
rect 30322 41694 30334 41746
rect 33618 41694 33630 41746
rect 33682 41743 33694 41746
rect 34290 41743 34302 41746
rect 33682 41697 34302 41743
rect 33682 41694 33694 41697
rect 34290 41694 34302 41697
rect 34354 41694 34366 41746
rect 8206 41682 8258 41694
rect 22318 41682 22370 41694
rect 46174 41682 46226 41694
rect 47070 41746 47122 41758
rect 47070 41682 47122 41694
rect 1344 41578 58576 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 58576 41578
rect 1344 41492 58576 41526
rect 21422 41410 21474 41422
rect 17154 41358 17166 41410
rect 17218 41358 17230 41410
rect 21422 41346 21474 41358
rect 26014 41410 26066 41422
rect 26014 41346 26066 41358
rect 37550 41410 37602 41422
rect 37550 41346 37602 41358
rect 42030 41410 42082 41422
rect 42030 41346 42082 41358
rect 47294 41410 47346 41422
rect 47294 41346 47346 41358
rect 1710 41298 1762 41310
rect 20862 41298 20914 41310
rect 8530 41246 8542 41298
rect 8594 41246 8606 41298
rect 11666 41246 11678 41298
rect 11730 41246 11742 41298
rect 18834 41246 18846 41298
rect 18898 41246 18910 41298
rect 1710 41234 1762 41246
rect 20862 41234 20914 41246
rect 22542 41298 22594 41310
rect 23438 41298 23490 41310
rect 22754 41246 22766 41298
rect 22818 41246 22830 41298
rect 22542 41234 22594 41246
rect 23438 41234 23490 41246
rect 24222 41298 24274 41310
rect 24222 41234 24274 41246
rect 27806 41298 27858 41310
rect 27806 41234 27858 41246
rect 30046 41298 30098 41310
rect 34638 41298 34690 41310
rect 34066 41246 34078 41298
rect 34130 41246 34142 41298
rect 30046 41234 30098 41246
rect 34638 41234 34690 41246
rect 40462 41298 40514 41310
rect 48078 41298 48130 41310
rect 42578 41246 42590 41298
rect 42642 41246 42654 41298
rect 46610 41246 46622 41298
rect 46674 41246 46686 41298
rect 40462 41234 40514 41246
rect 48078 41234 48130 41246
rect 49086 41298 49138 41310
rect 49086 41234 49138 41246
rect 52894 41298 52946 41310
rect 52894 41234 52946 41246
rect 57934 41298 57986 41310
rect 57934 41234 57986 41246
rect 17950 41186 18002 41198
rect 21534 41186 21586 41198
rect 7074 41134 7086 41186
rect 7138 41134 7150 41186
rect 8306 41134 8318 41186
rect 8370 41134 8382 41186
rect 8978 41134 8990 41186
rect 9042 41134 9054 41186
rect 10546 41134 10558 41186
rect 10610 41134 10622 41186
rect 11442 41134 11454 41186
rect 11506 41134 11518 41186
rect 12674 41134 12686 41186
rect 12738 41134 12750 41186
rect 13458 41134 13470 41186
rect 13522 41134 13534 41186
rect 14354 41134 14366 41186
rect 14418 41134 14430 41186
rect 14802 41134 14814 41186
rect 14866 41134 14878 41186
rect 16034 41134 16046 41186
rect 16098 41134 16110 41186
rect 17154 41134 17166 41186
rect 17218 41134 17230 41186
rect 17378 41134 17390 41186
rect 17442 41134 17454 41186
rect 18162 41134 18174 41186
rect 18226 41134 18238 41186
rect 18946 41134 18958 41186
rect 19010 41134 19022 41186
rect 17950 41122 18002 41134
rect 21534 41122 21586 41134
rect 22318 41186 22370 41198
rect 27022 41186 27074 41198
rect 33630 41186 33682 41198
rect 22866 41134 22878 41186
rect 22930 41134 22942 41186
rect 24546 41134 24558 41186
rect 24610 41134 24622 41186
rect 25442 41134 25454 41186
rect 25506 41134 25518 41186
rect 29586 41134 29598 41186
rect 29650 41134 29662 41186
rect 30594 41134 30606 41186
rect 30658 41134 30670 41186
rect 31490 41134 31502 41186
rect 31554 41134 31566 41186
rect 32610 41134 32622 41186
rect 32674 41134 32686 41186
rect 22318 41122 22370 41134
rect 27022 41122 27074 41134
rect 33630 41122 33682 41134
rect 34414 41186 34466 41198
rect 34414 41122 34466 41134
rect 34750 41186 34802 41198
rect 34750 41122 34802 41134
rect 35086 41186 35138 41198
rect 35086 41122 35138 41134
rect 37214 41186 37266 41198
rect 37214 41122 37266 41134
rect 38782 41186 38834 41198
rect 39678 41186 39730 41198
rect 41694 41186 41746 41198
rect 47518 41186 47570 41198
rect 39218 41134 39230 41186
rect 39282 41134 39294 41186
rect 40898 41134 40910 41186
rect 40962 41134 40974 41186
rect 42914 41134 42926 41186
rect 42978 41134 42990 41186
rect 45602 41134 45614 41186
rect 45666 41134 45678 41186
rect 46386 41134 46398 41186
rect 46450 41134 46462 41186
rect 38782 41122 38834 41134
rect 39678 41122 39730 41134
rect 41694 41122 41746 41134
rect 47518 41122 47570 41134
rect 47854 41186 47906 41198
rect 47854 41122 47906 41134
rect 48638 41186 48690 41198
rect 54574 41186 54626 41198
rect 52658 41134 52670 41186
rect 52722 41134 52734 41186
rect 56018 41134 56030 41186
rect 56082 41134 56094 41186
rect 48638 41122 48690 41134
rect 54574 41122 54626 41134
rect 21422 41074 21474 41086
rect 7298 41022 7310 41074
rect 7362 41022 7374 41074
rect 9202 41022 9214 41074
rect 9266 41022 9278 41074
rect 9650 41022 9662 41074
rect 9714 41022 9726 41074
rect 14242 41022 14254 41074
rect 14306 41022 14318 41074
rect 19618 41022 19630 41074
rect 19682 41022 19694 41074
rect 21422 41010 21474 41022
rect 26238 41074 26290 41086
rect 26238 41010 26290 41022
rect 26686 41074 26738 41086
rect 26686 41010 26738 41022
rect 28702 41074 28754 41086
rect 36990 41074 37042 41086
rect 43486 41074 43538 41086
rect 51326 41074 51378 41086
rect 30818 41022 30830 41074
rect 30882 41022 30894 41074
rect 31154 41022 31166 41074
rect 31218 41022 31230 41074
rect 41122 41022 41134 41074
rect 41186 41022 41198 41074
rect 46722 41022 46734 41074
rect 46786 41022 46798 41074
rect 28702 41010 28754 41022
rect 36990 41010 37042 41022
rect 43486 41010 43538 41022
rect 51326 41010 51378 41022
rect 51550 41074 51602 41086
rect 51550 41010 51602 41022
rect 51774 41074 51826 41086
rect 51774 41010 51826 41022
rect 51886 41074 51938 41086
rect 51886 41010 51938 41022
rect 53006 41074 53058 41086
rect 53006 41010 53058 41022
rect 53342 41074 53394 41086
rect 53342 41010 53394 41022
rect 54350 41074 54402 41086
rect 54350 41010 54402 41022
rect 54462 41074 54514 41086
rect 54462 41010 54514 41022
rect 20078 40962 20130 40974
rect 25678 40962 25730 40974
rect 24770 40910 24782 40962
rect 24834 40910 24846 40962
rect 20078 40898 20130 40910
rect 25678 40898 25730 40910
rect 26126 40962 26178 40974
rect 26126 40898 26178 40910
rect 26798 40962 26850 40974
rect 26798 40898 26850 40910
rect 27358 40962 27410 40974
rect 36542 40962 36594 40974
rect 31490 40910 31502 40962
rect 31554 40910 31566 40962
rect 27358 40898 27410 40910
rect 36542 40898 36594 40910
rect 48190 40962 48242 40974
rect 48190 40898 48242 40910
rect 53454 40962 53506 40974
rect 55010 40910 55022 40962
rect 55074 40910 55086 40962
rect 53454 40898 53506 40910
rect 1344 40794 58576 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 58576 40794
rect 1344 40708 58576 40742
rect 7198 40626 7250 40638
rect 7198 40562 7250 40574
rect 8878 40626 8930 40638
rect 12798 40626 12850 40638
rect 9874 40574 9886 40626
rect 9938 40574 9950 40626
rect 8878 40562 8930 40574
rect 12798 40562 12850 40574
rect 16270 40626 16322 40638
rect 16270 40562 16322 40574
rect 16382 40626 16434 40638
rect 16382 40562 16434 40574
rect 16494 40626 16546 40638
rect 16494 40562 16546 40574
rect 20750 40626 20802 40638
rect 22990 40626 23042 40638
rect 22194 40574 22206 40626
rect 22258 40574 22270 40626
rect 22418 40574 22430 40626
rect 22482 40574 22494 40626
rect 20750 40562 20802 40574
rect 22990 40562 23042 40574
rect 26574 40626 26626 40638
rect 29710 40626 29762 40638
rect 28690 40574 28702 40626
rect 28754 40574 28766 40626
rect 26574 40562 26626 40574
rect 29710 40562 29762 40574
rect 30270 40626 30322 40638
rect 30270 40562 30322 40574
rect 30606 40626 30658 40638
rect 30606 40562 30658 40574
rect 30830 40626 30882 40638
rect 30830 40562 30882 40574
rect 32062 40626 32114 40638
rect 32062 40562 32114 40574
rect 34190 40626 34242 40638
rect 34190 40562 34242 40574
rect 34862 40626 34914 40638
rect 34862 40562 34914 40574
rect 41694 40626 41746 40638
rect 41694 40562 41746 40574
rect 41806 40626 41858 40638
rect 41806 40562 41858 40574
rect 41918 40626 41970 40638
rect 41918 40562 41970 40574
rect 42142 40626 42194 40638
rect 42142 40562 42194 40574
rect 49982 40626 50034 40638
rect 49982 40562 50034 40574
rect 50990 40626 51042 40638
rect 53454 40626 53506 40638
rect 52098 40574 52110 40626
rect 52162 40574 52174 40626
rect 50990 40562 51042 40574
rect 53454 40562 53506 40574
rect 53678 40626 53730 40638
rect 55234 40574 55246 40626
rect 55298 40574 55310 40626
rect 53678 40562 53730 40574
rect 27134 40514 27186 40526
rect 7522 40462 7534 40514
rect 7586 40462 7598 40514
rect 10210 40462 10222 40514
rect 10274 40462 10286 40514
rect 21186 40462 21198 40514
rect 21250 40462 21262 40514
rect 27134 40450 27186 40462
rect 27358 40514 27410 40526
rect 31278 40514 31330 40526
rect 27682 40462 27694 40514
rect 27746 40462 27758 40514
rect 28354 40462 28366 40514
rect 28418 40462 28430 40514
rect 28578 40462 28590 40514
rect 28642 40462 28654 40514
rect 27358 40450 27410 40462
rect 31278 40450 31330 40462
rect 31838 40514 31890 40526
rect 31838 40450 31890 40462
rect 34974 40514 35026 40526
rect 34974 40450 35026 40462
rect 45838 40514 45890 40526
rect 45838 40450 45890 40462
rect 49422 40514 49474 40526
rect 49422 40450 49474 40462
rect 50542 40514 50594 40526
rect 50542 40450 50594 40462
rect 51662 40514 51714 40526
rect 51662 40450 51714 40462
rect 53342 40514 53394 40526
rect 56590 40514 56642 40526
rect 54450 40462 54462 40514
rect 54514 40462 54526 40514
rect 53342 40450 53394 40462
rect 56590 40450 56642 40462
rect 16942 40402 16994 40414
rect 23774 40402 23826 40414
rect 10098 40350 10110 40402
rect 10162 40350 10174 40402
rect 11330 40350 11342 40402
rect 11394 40350 11406 40402
rect 12002 40350 12014 40402
rect 12066 40350 12078 40402
rect 12674 40350 12686 40402
rect 12738 40350 12750 40402
rect 13682 40350 13694 40402
rect 13746 40350 13758 40402
rect 14802 40350 14814 40402
rect 14866 40350 14878 40402
rect 15810 40350 15822 40402
rect 15874 40350 15886 40402
rect 17826 40350 17838 40402
rect 17890 40350 17902 40402
rect 19282 40350 19294 40402
rect 19346 40350 19358 40402
rect 21634 40350 21646 40402
rect 21698 40350 21710 40402
rect 22082 40350 22094 40402
rect 22146 40350 22158 40402
rect 16942 40338 16994 40350
rect 23774 40338 23826 40350
rect 24334 40402 24386 40414
rect 25678 40402 25730 40414
rect 30494 40402 30546 40414
rect 25330 40350 25342 40402
rect 25394 40350 25406 40402
rect 25778 40350 25790 40402
rect 25842 40350 25854 40402
rect 28018 40350 28030 40402
rect 28082 40350 28094 40402
rect 24334 40338 24386 40350
rect 25678 40338 25730 40350
rect 30494 40338 30546 40350
rect 31166 40402 31218 40414
rect 31166 40338 31218 40350
rect 31502 40402 31554 40414
rect 31502 40338 31554 40350
rect 31726 40402 31778 40414
rect 31726 40338 31778 40350
rect 32174 40402 32226 40414
rect 32174 40338 32226 40350
rect 35086 40402 35138 40414
rect 35086 40338 35138 40350
rect 35198 40402 35250 40414
rect 46734 40402 46786 40414
rect 35410 40350 35422 40402
rect 35474 40350 35486 40402
rect 38322 40350 38334 40402
rect 38386 40350 38398 40402
rect 45266 40350 45278 40402
rect 45330 40350 45342 40402
rect 46274 40350 46286 40402
rect 46338 40350 46350 40402
rect 35198 40338 35250 40350
rect 46734 40338 46786 40350
rect 48862 40402 48914 40414
rect 48862 40338 48914 40350
rect 49310 40402 49362 40414
rect 49310 40338 49362 40350
rect 49534 40402 49586 40414
rect 51550 40402 51602 40414
rect 56926 40402 56978 40414
rect 50754 40350 50766 40402
rect 50818 40350 50830 40402
rect 51314 40350 51326 40402
rect 51378 40350 51390 40402
rect 54562 40350 54574 40402
rect 54626 40350 54638 40402
rect 55122 40350 55134 40402
rect 55186 40350 55198 40402
rect 49534 40338 49586 40350
rect 51550 40338 51602 40350
rect 56926 40338 56978 40350
rect 8206 40290 8258 40302
rect 44494 40290 44546 40302
rect 56814 40290 56866 40302
rect 17378 40238 17390 40290
rect 17442 40238 17454 40290
rect 19730 40238 19742 40290
rect 19794 40238 19806 40290
rect 37986 40238 37998 40290
rect 38050 40238 38062 40290
rect 44930 40238 44942 40290
rect 44994 40238 45006 40290
rect 8206 40226 8258 40238
rect 44494 40226 44546 40238
rect 56814 40226 56866 40238
rect 8094 40178 8146 40190
rect 8094 40114 8146 40126
rect 8430 40178 8482 40190
rect 51102 40178 51154 40190
rect 14914 40126 14926 40178
rect 14978 40126 14990 40178
rect 38658 40126 38670 40178
rect 38722 40126 38734 40178
rect 8430 40114 8482 40126
rect 51102 40114 51154 40126
rect 1344 40010 58576 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 58576 40010
rect 1344 39924 58576 39958
rect 9774 39842 9826 39854
rect 9774 39778 9826 39790
rect 11342 39842 11394 39854
rect 11342 39778 11394 39790
rect 22654 39842 22706 39854
rect 22654 39778 22706 39790
rect 23214 39842 23266 39854
rect 23214 39778 23266 39790
rect 23438 39842 23490 39854
rect 23438 39778 23490 39790
rect 29374 39842 29426 39854
rect 29374 39778 29426 39790
rect 29598 39842 29650 39854
rect 37998 39842 38050 39854
rect 37314 39790 37326 39842
rect 37378 39839 37390 39842
rect 37538 39839 37550 39842
rect 37378 39793 37550 39839
rect 37378 39790 37390 39793
rect 37538 39790 37550 39793
rect 37602 39790 37614 39842
rect 29598 39778 29650 39790
rect 37998 39778 38050 39790
rect 38334 39842 38386 39854
rect 38334 39778 38386 39790
rect 42366 39842 42418 39854
rect 42366 39778 42418 39790
rect 49086 39842 49138 39854
rect 54126 39842 54178 39854
rect 49746 39790 49758 39842
rect 49810 39790 49822 39842
rect 49086 39778 49138 39790
rect 54126 39778 54178 39790
rect 20750 39730 20802 39742
rect 12786 39678 12798 39730
rect 12850 39678 12862 39730
rect 19170 39678 19182 39730
rect 19234 39678 19246 39730
rect 20750 39666 20802 39678
rect 22430 39730 22482 39742
rect 22430 39666 22482 39678
rect 23102 39730 23154 39742
rect 23102 39666 23154 39678
rect 24222 39730 24274 39742
rect 24222 39666 24274 39678
rect 25006 39730 25058 39742
rect 25006 39666 25058 39678
rect 26014 39730 26066 39742
rect 31726 39730 31778 39742
rect 35870 39730 35922 39742
rect 28018 39678 28030 39730
rect 28082 39678 28094 39730
rect 33506 39678 33518 39730
rect 33570 39678 33582 39730
rect 26014 39666 26066 39678
rect 31726 39666 31778 39678
rect 35870 39666 35922 39678
rect 49198 39730 49250 39742
rect 57934 39730 57986 39742
rect 49858 39678 49870 39730
rect 49922 39678 49934 39730
rect 49198 39666 49250 39678
rect 57934 39666 57986 39678
rect 13470 39618 13522 39630
rect 6626 39566 6638 39618
rect 6690 39566 6702 39618
rect 7298 39566 7310 39618
rect 7362 39566 7374 39618
rect 7970 39566 7982 39618
rect 8034 39566 8046 39618
rect 8642 39566 8654 39618
rect 8706 39566 8718 39618
rect 9202 39566 9214 39618
rect 9266 39566 9278 39618
rect 9986 39566 9998 39618
rect 10050 39566 10062 39618
rect 10658 39566 10670 39618
rect 10722 39566 10734 39618
rect 11890 39566 11902 39618
rect 11954 39566 11966 39618
rect 13470 39554 13522 39566
rect 14030 39618 14082 39630
rect 21646 39618 21698 39630
rect 14690 39566 14702 39618
rect 14754 39566 14766 39618
rect 15362 39566 15374 39618
rect 15426 39566 15438 39618
rect 16594 39566 16606 39618
rect 16658 39566 16670 39618
rect 16930 39566 16942 39618
rect 16994 39566 17006 39618
rect 19282 39566 19294 39618
rect 19346 39566 19358 39618
rect 21298 39566 21310 39618
rect 21362 39566 21374 39618
rect 14030 39554 14082 39566
rect 21646 39554 21698 39566
rect 21982 39618 22034 39630
rect 21982 39554 22034 39566
rect 22094 39618 22146 39630
rect 22094 39554 22146 39566
rect 22206 39618 22258 39630
rect 24446 39618 24498 39630
rect 23650 39566 23662 39618
rect 23714 39566 23726 39618
rect 22206 39554 22258 39566
rect 24446 39554 24498 39566
rect 27694 39618 27746 39630
rect 34862 39618 34914 39630
rect 27906 39566 27918 39618
rect 27970 39566 27982 39618
rect 29138 39566 29150 39618
rect 29202 39566 29214 39618
rect 32050 39566 32062 39618
rect 32114 39566 32126 39618
rect 34290 39566 34302 39618
rect 34354 39566 34366 39618
rect 27694 39554 27746 39566
rect 34862 39554 34914 39566
rect 35422 39618 35474 39630
rect 35422 39554 35474 39566
rect 37774 39618 37826 39630
rect 37774 39554 37826 39566
rect 39566 39618 39618 39630
rect 39566 39554 39618 39566
rect 42142 39618 42194 39630
rect 42142 39554 42194 39566
rect 45166 39618 45218 39630
rect 48414 39618 48466 39630
rect 45826 39566 45838 39618
rect 45890 39566 45902 39618
rect 46722 39566 46734 39618
rect 46786 39566 46798 39618
rect 45166 39554 45218 39566
rect 48414 39554 48466 39566
rect 48638 39618 48690 39630
rect 48638 39554 48690 39566
rect 51102 39618 51154 39630
rect 56018 39566 56030 39618
rect 56082 39566 56094 39618
rect 51102 39554 51154 39566
rect 25118 39506 25170 39518
rect 6850 39454 6862 39506
rect 6914 39454 6926 39506
rect 8194 39454 8206 39506
rect 8258 39454 8270 39506
rect 14578 39454 14590 39506
rect 14642 39454 14654 39506
rect 19730 39454 19742 39506
rect 19794 39454 19806 39506
rect 25118 39442 25170 39454
rect 29710 39506 29762 39518
rect 35758 39506 35810 39518
rect 48974 39506 49026 39518
rect 50990 39506 51042 39518
rect 32274 39454 32286 39506
rect 32338 39454 32350 39506
rect 45938 39454 45950 39506
rect 46002 39454 46014 39506
rect 49634 39454 49646 39506
rect 49698 39454 49710 39506
rect 29710 39442 29762 39454
rect 35758 39442 35810 39454
rect 48974 39442 49026 39454
rect 50990 39442 51042 39454
rect 54238 39506 54290 39518
rect 54238 39442 54290 39454
rect 1710 39394 1762 39406
rect 24894 39394 24946 39406
rect 7522 39342 7534 39394
rect 7586 39342 7598 39394
rect 15474 39342 15486 39394
rect 15538 39342 15550 39394
rect 1710 39330 1762 39342
rect 24894 39330 24946 39342
rect 28590 39394 28642 39406
rect 28590 39330 28642 39342
rect 35982 39394 36034 39406
rect 54126 39394 54178 39406
rect 39890 39342 39902 39394
rect 39954 39342 39966 39394
rect 42690 39342 42702 39394
rect 42754 39342 42766 39394
rect 44818 39342 44830 39394
rect 44882 39342 44894 39394
rect 46834 39342 46846 39394
rect 46898 39342 46910 39394
rect 35982 39330 36034 39342
rect 54126 39330 54178 39342
rect 1344 39226 58576 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 58576 39226
rect 1344 39140 58576 39174
rect 9550 39058 9602 39070
rect 9550 38994 9602 39006
rect 10782 39058 10834 39070
rect 10782 38994 10834 39006
rect 11678 39058 11730 39070
rect 11678 38994 11730 39006
rect 12574 39058 12626 39070
rect 12574 38994 12626 39006
rect 13470 39058 13522 39070
rect 13470 38994 13522 39006
rect 16270 39058 16322 39070
rect 19182 39058 19234 39070
rect 18386 39006 18398 39058
rect 18450 39006 18462 39058
rect 16270 38994 16322 39006
rect 19182 38994 19234 39006
rect 19518 39058 19570 39070
rect 19518 38994 19570 39006
rect 20750 39058 20802 39070
rect 20750 38994 20802 39006
rect 22206 39058 22258 39070
rect 22206 38994 22258 39006
rect 22430 39058 22482 39070
rect 22430 38994 22482 39006
rect 22654 39058 22706 39070
rect 22654 38994 22706 39006
rect 23998 39058 24050 39070
rect 23998 38994 24050 39006
rect 33406 39058 33458 39070
rect 33406 38994 33458 39006
rect 33854 39058 33906 39070
rect 33854 38994 33906 39006
rect 35198 39058 35250 39070
rect 47854 39058 47906 39070
rect 42578 39006 42590 39058
rect 42642 39006 42654 39058
rect 43586 39006 43598 39058
rect 43650 39006 43662 39058
rect 35198 38994 35250 39006
rect 47854 38994 47906 39006
rect 49646 39058 49698 39070
rect 49646 38994 49698 39006
rect 50094 39058 50146 39070
rect 50094 38994 50146 39006
rect 53230 39058 53282 39070
rect 53230 38994 53282 39006
rect 7646 38946 7698 38958
rect 7646 38882 7698 38894
rect 16830 38946 16882 38958
rect 20862 38946 20914 38958
rect 17826 38894 17838 38946
rect 17890 38894 17902 38946
rect 16830 38882 16882 38894
rect 20862 38882 20914 38894
rect 22878 38946 22930 38958
rect 35758 38946 35810 38958
rect 43038 38946 43090 38958
rect 50542 38946 50594 38958
rect 28466 38894 28478 38946
rect 28530 38894 28542 38946
rect 34850 38894 34862 38946
rect 34914 38894 34926 38946
rect 41794 38894 41806 38946
rect 41858 38894 41870 38946
rect 45602 38894 45614 38946
rect 45666 38894 45678 38946
rect 46274 38894 46286 38946
rect 46338 38894 46350 38946
rect 22878 38882 22930 38894
rect 35758 38882 35810 38894
rect 43038 38882 43090 38894
rect 50542 38882 50594 38894
rect 54798 38946 54850 38958
rect 54798 38882 54850 38894
rect 11342 38834 11394 38846
rect 11342 38770 11394 38782
rect 12238 38834 12290 38846
rect 12238 38770 12290 38782
rect 14030 38834 14082 38846
rect 14030 38770 14082 38782
rect 14814 38834 14866 38846
rect 14814 38770 14866 38782
rect 15262 38834 15314 38846
rect 22990 38834 23042 38846
rect 29262 38834 29314 38846
rect 31726 38834 31778 38846
rect 17938 38782 17950 38834
rect 18002 38782 18014 38834
rect 18274 38782 18286 38834
rect 18338 38782 18350 38834
rect 21858 38782 21870 38834
rect 21922 38782 21934 38834
rect 24098 38782 24110 38834
rect 24162 38782 24174 38834
rect 27794 38782 27806 38834
rect 27858 38782 27870 38834
rect 29474 38782 29486 38834
rect 29538 38782 29550 38834
rect 15262 38770 15314 38782
rect 22990 38770 23042 38782
rect 29262 38770 29314 38782
rect 31726 38770 31778 38782
rect 31950 38834 32002 38846
rect 31950 38770 32002 38782
rect 32286 38834 32338 38846
rect 32286 38770 32338 38782
rect 35534 38834 35586 38846
rect 35534 38770 35586 38782
rect 36094 38834 36146 38846
rect 43262 38834 43314 38846
rect 45054 38834 45106 38846
rect 38546 38782 38558 38834
rect 38610 38782 38622 38834
rect 42130 38782 42142 38834
rect 42194 38782 42206 38834
rect 42466 38782 42478 38834
rect 42530 38782 42542 38834
rect 44706 38782 44718 38834
rect 44770 38782 44782 38834
rect 36094 38770 36146 38782
rect 43262 38770 43314 38782
rect 45054 38770 45106 38782
rect 45166 38834 45218 38846
rect 48974 38834 49026 38846
rect 45938 38782 45950 38834
rect 46002 38782 46014 38834
rect 46386 38782 46398 38834
rect 46450 38782 46462 38834
rect 47282 38782 47294 38834
rect 47346 38782 47358 38834
rect 45166 38770 45218 38782
rect 48974 38770 49026 38782
rect 49198 38834 49250 38846
rect 49198 38770 49250 38782
rect 53118 38834 53170 38846
rect 53118 38770 53170 38782
rect 53454 38834 53506 38846
rect 54114 38782 54126 38834
rect 54178 38782 54190 38834
rect 53454 38770 53506 38782
rect 8430 38722 8482 38734
rect 13134 38722 13186 38734
rect 22318 38722 22370 38734
rect 32510 38722 32562 38734
rect 7858 38670 7870 38722
rect 7922 38670 7934 38722
rect 9986 38670 9998 38722
rect 10050 38670 10062 38722
rect 19954 38670 19966 38722
rect 20018 38670 20030 38722
rect 23986 38670 23998 38722
rect 24050 38670 24062 38722
rect 8430 38658 8482 38670
rect 13134 38658 13186 38670
rect 22318 38658 22370 38670
rect 32510 38658 32562 38670
rect 35982 38722 36034 38734
rect 39230 38722 39282 38734
rect 38322 38670 38334 38722
rect 38386 38670 38398 38722
rect 35982 38658 36034 38670
rect 39230 38658 39282 38670
rect 48750 38722 48802 38734
rect 54002 38670 54014 38722
rect 54066 38670 54078 38722
rect 48750 38658 48802 38670
rect 20638 38610 20690 38622
rect 32398 38610 32450 38622
rect 14578 38558 14590 38610
rect 14642 38558 14654 38610
rect 27682 38558 27694 38610
rect 27746 38558 27758 38610
rect 20638 38546 20690 38558
rect 32398 38546 32450 38558
rect 1344 38442 58576 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 58576 38442
rect 1344 38356 58576 38390
rect 14814 38274 14866 38286
rect 15138 38222 15150 38274
rect 15202 38222 15214 38274
rect 33282 38222 33294 38274
rect 33346 38222 33358 38274
rect 46050 38222 46062 38274
rect 46114 38222 46126 38274
rect 53218 38222 53230 38274
rect 53282 38222 53294 38274
rect 14814 38210 14866 38222
rect 14590 38162 14642 38174
rect 14590 38098 14642 38110
rect 16158 38162 16210 38174
rect 16158 38098 16210 38110
rect 17054 38162 17106 38174
rect 17054 38098 17106 38110
rect 19294 38162 19346 38174
rect 19294 38098 19346 38110
rect 24558 38162 24610 38174
rect 30158 38162 30210 38174
rect 34190 38162 34242 38174
rect 51886 38162 51938 38174
rect 27906 38110 27918 38162
rect 27970 38110 27982 38162
rect 32162 38110 32174 38162
rect 32226 38110 32238 38162
rect 35746 38110 35758 38162
rect 35810 38110 35822 38162
rect 43362 38110 43374 38162
rect 43426 38110 43438 38162
rect 45266 38110 45278 38162
rect 45330 38110 45342 38162
rect 51426 38110 51438 38162
rect 51490 38110 51502 38162
rect 53554 38110 53566 38162
rect 53618 38110 53630 38162
rect 57698 38110 57710 38162
rect 57762 38110 57774 38162
rect 24558 38098 24610 38110
rect 30158 38098 30210 38110
rect 34190 38098 34242 38110
rect 51886 38098 51938 38110
rect 14030 38050 14082 38062
rect 17838 38050 17890 38062
rect 16594 37998 16606 38050
rect 16658 37998 16670 38050
rect 14030 37986 14082 37998
rect 17838 37986 17890 37998
rect 18734 38050 18786 38062
rect 18734 37986 18786 37998
rect 20750 38050 20802 38062
rect 20750 37986 20802 37998
rect 21870 38050 21922 38062
rect 21870 37986 21922 37998
rect 23438 38050 23490 38062
rect 23438 37986 23490 37998
rect 24782 38050 24834 38062
rect 24782 37986 24834 37998
rect 25230 38050 25282 38062
rect 25230 37986 25282 37998
rect 25454 38050 25506 38062
rect 25454 37986 25506 37998
rect 26238 38050 26290 38062
rect 29038 38050 29090 38062
rect 26562 37998 26574 38050
rect 26626 37998 26638 38050
rect 27122 37998 27134 38050
rect 27186 37998 27198 38050
rect 28578 37998 28590 38050
rect 28642 37998 28654 38050
rect 26238 37986 26290 37998
rect 29038 37986 29090 37998
rect 29262 38050 29314 38062
rect 29262 37986 29314 37998
rect 29374 38050 29426 38062
rect 29374 37986 29426 37998
rect 31166 38050 31218 38062
rect 32846 38050 32898 38062
rect 37550 38050 37602 38062
rect 31714 37998 31726 38050
rect 31778 37998 31790 38050
rect 32050 37998 32062 38050
rect 32114 37998 32126 38050
rect 33058 37998 33070 38050
rect 33122 37998 33134 38050
rect 34514 37998 34526 38050
rect 34578 37998 34590 38050
rect 34850 37998 34862 38050
rect 34914 37998 34926 38050
rect 35858 37998 35870 38050
rect 35922 37998 35934 38050
rect 31166 37986 31218 37998
rect 32846 37986 32898 37998
rect 37550 37986 37602 37998
rect 37886 38050 37938 38062
rect 37886 37986 37938 37998
rect 38110 38050 38162 38062
rect 43262 38050 43314 38062
rect 53454 38050 53506 38062
rect 42466 37998 42478 38050
rect 42530 37998 42542 38050
rect 43474 37998 43486 38050
rect 43538 37998 43550 38050
rect 45378 37998 45390 38050
rect 45442 37998 45454 38050
rect 51202 37998 51214 38050
rect 51266 37998 51278 38050
rect 38110 37986 38162 37998
rect 43262 37986 43314 37998
rect 53454 37986 53506 37998
rect 54350 38050 54402 38062
rect 54562 37998 54574 38050
rect 54626 37998 54638 38050
rect 55794 37998 55806 38050
rect 55858 37998 55870 38050
rect 54350 37986 54402 37998
rect 10222 37938 10274 37950
rect 10222 37874 10274 37886
rect 18398 37938 18450 37950
rect 18398 37874 18450 37886
rect 23998 37938 24050 37950
rect 29710 37938 29762 37950
rect 42254 37938 42306 37950
rect 28130 37886 28142 37938
rect 28194 37886 28206 37938
rect 34962 37886 34974 37938
rect 35026 37886 35038 37938
rect 35634 37886 35646 37938
rect 35698 37886 35710 37938
rect 23998 37874 24050 37886
rect 29710 37874 29762 37886
rect 42254 37874 42306 37886
rect 55246 37938 55298 37950
rect 55246 37874 55298 37886
rect 13470 37826 13522 37838
rect 10546 37774 10558 37826
rect 10610 37774 10622 37826
rect 13470 37762 13522 37774
rect 15598 37826 15650 37838
rect 15598 37762 15650 37774
rect 19742 37826 19794 37838
rect 19742 37762 19794 37774
rect 20190 37826 20242 37838
rect 20190 37762 20242 37774
rect 21310 37826 21362 37838
rect 21310 37762 21362 37774
rect 25342 37826 25394 37838
rect 25342 37762 25394 37774
rect 26014 37826 26066 37838
rect 26014 37762 26066 37774
rect 26798 37826 26850 37838
rect 26798 37762 26850 37774
rect 26910 37826 26962 37838
rect 26910 37762 26962 37774
rect 27358 37826 27410 37838
rect 27358 37762 27410 37774
rect 34302 37826 34354 37838
rect 34302 37762 34354 37774
rect 37886 37826 37938 37838
rect 37886 37762 37938 37774
rect 1344 37658 58576 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 58576 37658
rect 1344 37572 58576 37606
rect 6974 37490 7026 37502
rect 6974 37426 7026 37438
rect 7646 37490 7698 37502
rect 17614 37490 17666 37502
rect 8642 37438 8654 37490
rect 8706 37438 8718 37490
rect 15922 37438 15934 37490
rect 15986 37438 15998 37490
rect 7646 37426 7698 37438
rect 17614 37426 17666 37438
rect 18734 37490 18786 37502
rect 23550 37490 23602 37502
rect 19058 37438 19070 37490
rect 19122 37438 19134 37490
rect 22082 37438 22094 37490
rect 22146 37438 22158 37490
rect 18734 37426 18786 37438
rect 23550 37426 23602 37438
rect 23998 37490 24050 37502
rect 23998 37426 24050 37438
rect 24334 37490 24386 37502
rect 24334 37426 24386 37438
rect 27470 37490 27522 37502
rect 27470 37426 27522 37438
rect 28254 37490 28306 37502
rect 28254 37426 28306 37438
rect 33406 37490 33458 37502
rect 41358 37490 41410 37502
rect 37650 37438 37662 37490
rect 37714 37438 37726 37490
rect 40338 37438 40350 37490
rect 40402 37438 40414 37490
rect 33406 37426 33458 37438
rect 41358 37426 41410 37438
rect 50542 37490 50594 37502
rect 50542 37426 50594 37438
rect 50654 37490 50706 37502
rect 50654 37426 50706 37438
rect 54350 37490 54402 37502
rect 54350 37426 54402 37438
rect 56030 37490 56082 37502
rect 56030 37426 56082 37438
rect 1710 37378 1762 37390
rect 1710 37314 1762 37326
rect 14030 37378 14082 37390
rect 14030 37314 14082 37326
rect 15150 37378 15202 37390
rect 24222 37378 24274 37390
rect 19618 37326 19630 37378
rect 19682 37326 19694 37378
rect 15150 37314 15202 37326
rect 24222 37314 24274 37326
rect 29710 37378 29762 37390
rect 29710 37314 29762 37326
rect 30718 37378 30770 37390
rect 37214 37378 37266 37390
rect 39342 37378 39394 37390
rect 32162 37326 32174 37378
rect 32226 37326 32238 37378
rect 33058 37326 33070 37378
rect 33122 37326 33134 37378
rect 34066 37326 34078 37378
rect 34130 37326 34142 37378
rect 38434 37326 38446 37378
rect 38498 37326 38510 37378
rect 30718 37314 30770 37326
rect 37214 37314 37266 37326
rect 39342 37314 39394 37326
rect 44270 37378 44322 37390
rect 44270 37314 44322 37326
rect 49758 37378 49810 37390
rect 49758 37314 49810 37326
rect 51662 37378 51714 37390
rect 51662 37314 51714 37326
rect 54574 37378 54626 37390
rect 54574 37314 54626 37326
rect 54798 37378 54850 37390
rect 54798 37314 54850 37326
rect 55694 37378 55746 37390
rect 55694 37314 55746 37326
rect 10670 37266 10722 37278
rect 13134 37266 13186 37278
rect 15374 37266 15426 37278
rect 7186 37214 7198 37266
rect 7250 37214 7262 37266
rect 8866 37214 8878 37266
rect 8930 37214 8942 37266
rect 9650 37214 9662 37266
rect 9714 37214 9726 37266
rect 11106 37214 11118 37266
rect 11170 37214 11182 37266
rect 13570 37214 13582 37266
rect 13634 37214 13646 37266
rect 10670 37202 10722 37214
rect 13134 37202 13186 37214
rect 15374 37202 15426 37214
rect 15598 37266 15650 37278
rect 20526 37266 20578 37278
rect 24558 37266 24610 37278
rect 18274 37214 18286 37266
rect 18338 37214 18350 37266
rect 19842 37214 19854 37266
rect 19906 37214 19918 37266
rect 20738 37214 20750 37266
rect 20802 37214 20814 37266
rect 21858 37214 21870 37266
rect 21922 37214 21934 37266
rect 15598 37202 15650 37214
rect 20526 37202 20578 37214
rect 24558 37202 24610 37214
rect 26910 37266 26962 37278
rect 27582 37266 27634 37278
rect 27234 37214 27246 37266
rect 27298 37214 27310 37266
rect 26910 37202 26962 37214
rect 27582 37202 27634 37214
rect 27806 37266 27858 37278
rect 27806 37202 27858 37214
rect 28142 37266 28194 37278
rect 28142 37202 28194 37214
rect 28478 37266 28530 37278
rect 39006 37266 39058 37278
rect 28914 37214 28926 37266
rect 28978 37214 28990 37266
rect 30034 37214 30046 37266
rect 30098 37214 30110 37266
rect 30930 37214 30942 37266
rect 30994 37214 31006 37266
rect 32050 37214 32062 37266
rect 32114 37214 32126 37266
rect 33954 37214 33966 37266
rect 34018 37214 34030 37266
rect 36194 37214 36206 37266
rect 36258 37214 36270 37266
rect 38322 37214 38334 37266
rect 38386 37214 38398 37266
rect 28478 37202 28530 37214
rect 39006 37202 39058 37214
rect 39790 37266 39842 37278
rect 39790 37202 39842 37214
rect 41022 37266 41074 37278
rect 41022 37202 41074 37214
rect 41358 37266 41410 37278
rect 41358 37202 41410 37214
rect 41694 37266 41746 37278
rect 41694 37202 41746 37214
rect 42142 37266 42194 37278
rect 44158 37266 44210 37278
rect 42354 37214 42366 37266
rect 42418 37214 42430 37266
rect 42142 37202 42194 37214
rect 44158 37202 44210 37214
rect 44494 37266 44546 37278
rect 44494 37202 44546 37214
rect 44718 37266 44770 37278
rect 45726 37266 45778 37278
rect 50094 37266 50146 37278
rect 45266 37214 45278 37266
rect 45330 37214 45342 37266
rect 45938 37214 45950 37266
rect 46002 37214 46014 37266
rect 44718 37202 44770 37214
rect 45726 37202 45778 37214
rect 50094 37202 50146 37214
rect 50766 37266 50818 37278
rect 52894 37266 52946 37278
rect 51090 37214 51102 37266
rect 51154 37214 51166 37266
rect 50766 37202 50818 37214
rect 52894 37202 52946 37214
rect 54126 37266 54178 37278
rect 54126 37202 54178 37214
rect 8206 37154 8258 37166
rect 49870 37154 49922 37166
rect 9986 37102 9998 37154
rect 10050 37102 10062 37154
rect 12674 37102 12686 37154
rect 12738 37102 12750 37154
rect 17938 37102 17950 37154
rect 18002 37102 18014 37154
rect 20178 37102 20190 37154
rect 20242 37102 20254 37154
rect 29138 37102 29150 37154
rect 29202 37102 29214 37154
rect 30146 37102 30158 37154
rect 30210 37102 30222 37154
rect 31938 37102 31950 37154
rect 32002 37102 32014 37154
rect 46050 37102 46062 37154
rect 46114 37102 46126 37154
rect 8206 37090 8258 37102
rect 49870 37090 49922 37102
rect 53006 37154 53058 37166
rect 53006 37090 53058 37102
rect 2158 37042 2210 37054
rect 40014 37042 40066 37054
rect 21186 36990 21198 37042
rect 21250 36990 21262 37042
rect 2158 36978 2210 36990
rect 40014 36978 40066 36990
rect 42030 37042 42082 37054
rect 42030 36978 42082 36990
rect 1344 36874 58576 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 58576 36874
rect 1344 36788 58576 36822
rect 13918 36706 13970 36718
rect 13918 36642 13970 36654
rect 14590 36706 14642 36718
rect 14590 36642 14642 36654
rect 22094 36706 22146 36718
rect 22094 36642 22146 36654
rect 22318 36706 22370 36718
rect 22318 36642 22370 36654
rect 26238 36706 26290 36718
rect 26238 36642 26290 36654
rect 29486 36706 29538 36718
rect 29486 36642 29538 36654
rect 35086 36706 35138 36718
rect 35086 36642 35138 36654
rect 35422 36706 35474 36718
rect 35422 36642 35474 36654
rect 36094 36706 36146 36718
rect 54238 36706 54290 36718
rect 45938 36654 45950 36706
rect 46002 36654 46014 36706
rect 50978 36654 50990 36706
rect 51042 36654 51054 36706
rect 36094 36642 36146 36654
rect 54238 36642 54290 36654
rect 1934 36594 1986 36606
rect 1934 36530 1986 36542
rect 8990 36594 9042 36606
rect 11790 36594 11842 36606
rect 10994 36542 11006 36594
rect 11058 36542 11070 36594
rect 8990 36530 9042 36542
rect 11790 36530 11842 36542
rect 18846 36594 18898 36606
rect 20750 36594 20802 36606
rect 19394 36542 19406 36594
rect 19458 36542 19470 36594
rect 18846 36530 18898 36542
rect 20750 36530 20802 36542
rect 21534 36594 21586 36606
rect 30382 36594 30434 36606
rect 23538 36542 23550 36594
rect 23602 36542 23614 36594
rect 26562 36542 26574 36594
rect 26626 36542 26638 36594
rect 29250 36542 29262 36594
rect 29314 36542 29326 36594
rect 31042 36542 31054 36594
rect 31106 36542 31118 36594
rect 33506 36542 33518 36594
rect 33570 36542 33582 36594
rect 41794 36542 41806 36594
rect 41858 36542 41870 36594
rect 49298 36542 49310 36594
rect 49362 36542 49374 36594
rect 51426 36542 51438 36594
rect 51490 36542 51502 36594
rect 21534 36530 21586 36542
rect 30382 36530 30434 36542
rect 8430 36482 8482 36494
rect 12126 36482 12178 36494
rect 13470 36482 13522 36494
rect 4274 36430 4286 36482
rect 4338 36430 4350 36482
rect 9426 36430 9438 36482
rect 9490 36430 9502 36482
rect 9762 36430 9774 36482
rect 9826 36430 9838 36482
rect 12338 36430 12350 36482
rect 12402 36430 12414 36482
rect 8430 36418 8482 36430
rect 12126 36418 12178 36430
rect 13470 36418 13522 36430
rect 13694 36482 13746 36494
rect 13694 36418 13746 36430
rect 14142 36482 14194 36494
rect 20190 36482 20242 36494
rect 15474 36430 15486 36482
rect 15538 36430 15550 36482
rect 16370 36430 16382 36482
rect 16434 36430 16446 36482
rect 17154 36430 17166 36482
rect 17218 36430 17230 36482
rect 19730 36430 19742 36482
rect 19794 36430 19806 36482
rect 14142 36418 14194 36430
rect 20190 36418 20242 36430
rect 21870 36482 21922 36494
rect 27358 36482 27410 36494
rect 27918 36482 27970 36494
rect 22866 36430 22878 36482
rect 22930 36430 22942 36482
rect 23986 36430 23998 36482
rect 24050 36430 24062 36482
rect 24658 36430 24670 36482
rect 24722 36430 24734 36482
rect 25554 36430 25566 36482
rect 25618 36430 25630 36482
rect 27570 36430 27582 36482
rect 27634 36430 27646 36482
rect 21870 36418 21922 36430
rect 27358 36418 27410 36430
rect 27918 36418 27970 36430
rect 28254 36482 28306 36494
rect 33966 36482 34018 36494
rect 29138 36430 29150 36482
rect 29202 36430 29214 36482
rect 31378 36430 31390 36482
rect 31442 36430 31454 36482
rect 32386 36430 32398 36482
rect 32450 36430 32462 36482
rect 33282 36430 33294 36482
rect 33346 36430 33358 36482
rect 28254 36418 28306 36430
rect 33966 36418 34018 36430
rect 35198 36482 35250 36494
rect 51214 36482 51266 36494
rect 35634 36430 35646 36482
rect 35698 36430 35710 36482
rect 39330 36430 39342 36482
rect 39394 36430 39406 36482
rect 41570 36430 41582 36482
rect 41634 36430 41646 36482
rect 42242 36430 42254 36482
rect 42306 36430 42318 36482
rect 44818 36430 44830 36482
rect 44882 36430 44894 36482
rect 46050 36430 46062 36482
rect 46114 36430 46126 36482
rect 47058 36430 47070 36482
rect 47122 36430 47134 36482
rect 48514 36430 48526 36482
rect 48578 36430 48590 36482
rect 49522 36430 49534 36482
rect 49586 36430 49598 36482
rect 35198 36418 35250 36430
rect 51214 36418 51266 36430
rect 53566 36482 53618 36494
rect 53566 36418 53618 36430
rect 53902 36482 53954 36494
rect 55570 36430 55582 36482
rect 55634 36430 55646 36482
rect 53902 36418 53954 36430
rect 7534 36370 7586 36382
rect 7534 36306 7586 36318
rect 12910 36370 12962 36382
rect 22766 36370 22818 36382
rect 26462 36370 26514 36382
rect 15362 36318 15374 36370
rect 15426 36318 15438 36370
rect 15698 36318 15710 36370
rect 15762 36318 15774 36370
rect 16146 36318 16158 36370
rect 16210 36318 16222 36370
rect 18386 36318 18398 36370
rect 18450 36318 18462 36370
rect 24322 36318 24334 36370
rect 24386 36318 24398 36370
rect 24882 36318 24894 36370
rect 24946 36318 24958 36370
rect 12910 36306 12962 36318
rect 22766 36306 22818 36318
rect 26462 36306 26514 36318
rect 28142 36370 28194 36382
rect 28142 36306 28194 36318
rect 30718 36370 30770 36382
rect 30718 36306 30770 36318
rect 30942 36370 30994 36382
rect 34078 36370 34130 36382
rect 32610 36318 32622 36370
rect 32674 36318 32686 36370
rect 33170 36318 33182 36370
rect 33234 36318 33246 36370
rect 30942 36306 30994 36318
rect 34078 36306 34130 36318
rect 34414 36370 34466 36382
rect 34414 36306 34466 36318
rect 35982 36370 36034 36382
rect 35982 36306 36034 36318
rect 36094 36370 36146 36382
rect 36094 36306 36146 36318
rect 37998 36370 38050 36382
rect 53790 36370 53842 36382
rect 39106 36318 39118 36370
rect 39170 36318 39182 36370
rect 42578 36318 42590 36370
rect 42642 36318 42654 36370
rect 47282 36318 47294 36370
rect 47346 36318 47358 36370
rect 49186 36318 49198 36370
rect 49250 36318 49262 36370
rect 37998 36306 38050 36318
rect 53790 36306 53842 36318
rect 54350 36370 54402 36382
rect 54350 36306 54402 36318
rect 7870 36258 7922 36270
rect 17726 36258 17778 36270
rect 17042 36206 17054 36258
rect 17106 36206 17118 36258
rect 7870 36194 7922 36206
rect 17726 36194 17778 36206
rect 18062 36258 18114 36270
rect 27022 36258 27074 36270
rect 25666 36206 25678 36258
rect 25730 36206 25742 36258
rect 18062 36194 18114 36206
rect 27022 36194 27074 36206
rect 29934 36258 29986 36270
rect 29934 36194 29986 36206
rect 34190 36258 34242 36270
rect 34190 36194 34242 36206
rect 38110 36258 38162 36270
rect 38110 36194 38162 36206
rect 38334 36258 38386 36270
rect 56590 36258 56642 36270
rect 39554 36206 39566 36258
rect 39618 36206 39630 36258
rect 38334 36194 38386 36206
rect 56590 36194 56642 36206
rect 1344 36090 58576 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 58576 36090
rect 1344 36004 58576 36038
rect 17390 35922 17442 35934
rect 8194 35870 8206 35922
rect 8258 35870 8270 35922
rect 14242 35870 14254 35922
rect 14306 35870 14318 35922
rect 16258 35870 16270 35922
rect 16322 35870 16334 35922
rect 17390 35858 17442 35870
rect 19070 35922 19122 35934
rect 19070 35858 19122 35870
rect 19854 35922 19906 35934
rect 19854 35858 19906 35870
rect 21422 35922 21474 35934
rect 21422 35858 21474 35870
rect 24670 35922 24722 35934
rect 24670 35858 24722 35870
rect 25342 35922 25394 35934
rect 25342 35858 25394 35870
rect 27022 35922 27074 35934
rect 27022 35858 27074 35870
rect 27246 35922 27298 35934
rect 27246 35858 27298 35870
rect 28366 35922 28418 35934
rect 28366 35858 28418 35870
rect 28814 35922 28866 35934
rect 28814 35858 28866 35870
rect 29710 35922 29762 35934
rect 29710 35858 29762 35870
rect 30158 35922 30210 35934
rect 30158 35858 30210 35870
rect 34862 35922 34914 35934
rect 34862 35858 34914 35870
rect 36766 35922 36818 35934
rect 36766 35858 36818 35870
rect 41582 35922 41634 35934
rect 41582 35858 41634 35870
rect 42366 35922 42418 35934
rect 42366 35858 42418 35870
rect 10670 35810 10722 35822
rect 15710 35810 15762 35822
rect 13570 35758 13582 35810
rect 13634 35758 13646 35810
rect 14914 35758 14926 35810
rect 14978 35758 14990 35810
rect 10670 35746 10722 35758
rect 15710 35746 15762 35758
rect 22766 35810 22818 35822
rect 22766 35746 22818 35758
rect 25230 35810 25282 35822
rect 25230 35746 25282 35758
rect 26910 35810 26962 35822
rect 26910 35746 26962 35758
rect 29486 35810 29538 35822
rect 29486 35746 29538 35758
rect 30270 35810 30322 35822
rect 30270 35746 30322 35758
rect 36206 35810 36258 35822
rect 36206 35746 36258 35758
rect 37438 35810 37490 35822
rect 41246 35810 41298 35822
rect 39442 35758 39454 35810
rect 39506 35758 39518 35810
rect 37438 35746 37490 35758
rect 41246 35746 41298 35758
rect 41358 35810 41410 35822
rect 48078 35810 48130 35822
rect 43026 35758 43038 35810
rect 43090 35758 43102 35810
rect 41358 35746 41410 35758
rect 48078 35746 48130 35758
rect 49758 35810 49810 35822
rect 49758 35746 49810 35758
rect 6862 35698 6914 35710
rect 4274 35646 4286 35698
rect 4338 35646 4350 35698
rect 6862 35634 6914 35646
rect 7422 35698 7474 35710
rect 11118 35698 11170 35710
rect 8418 35646 8430 35698
rect 8482 35646 8494 35698
rect 9986 35646 9998 35698
rect 10050 35646 10062 35698
rect 7422 35634 7474 35646
rect 11118 35634 11170 35646
rect 11678 35698 11730 35710
rect 11678 35634 11730 35646
rect 12014 35698 12066 35710
rect 15934 35698 15986 35710
rect 13234 35646 13246 35698
rect 13298 35646 13310 35698
rect 14130 35646 14142 35698
rect 14194 35646 14206 35698
rect 14802 35646 14814 35698
rect 14866 35646 14878 35698
rect 12014 35634 12066 35646
rect 15934 35634 15986 35646
rect 20414 35698 20466 35710
rect 20414 35634 20466 35646
rect 25566 35698 25618 35710
rect 25566 35634 25618 35646
rect 29374 35698 29426 35710
rect 29374 35634 29426 35646
rect 29822 35698 29874 35710
rect 29822 35634 29874 35646
rect 30382 35698 30434 35710
rect 35758 35698 35810 35710
rect 33170 35646 33182 35698
rect 33234 35646 33246 35698
rect 33618 35646 33630 35698
rect 33682 35646 33694 35698
rect 34514 35646 34526 35698
rect 34578 35646 34590 35698
rect 35298 35646 35310 35698
rect 35362 35646 35374 35698
rect 30382 35634 30434 35646
rect 35758 35634 35810 35646
rect 37214 35698 37266 35710
rect 37214 35634 37266 35646
rect 37550 35698 37602 35710
rect 47182 35698 47234 35710
rect 52558 35698 52610 35710
rect 38322 35646 38334 35698
rect 38386 35646 38398 35698
rect 38770 35646 38782 35698
rect 38834 35646 38846 35698
rect 42802 35646 42814 35698
rect 42866 35646 42878 35698
rect 45714 35646 45726 35698
rect 45778 35646 45790 35698
rect 46274 35646 46286 35698
rect 46338 35646 46350 35698
rect 47394 35646 47406 35698
rect 47458 35646 47470 35698
rect 49074 35646 49086 35698
rect 49138 35646 49150 35698
rect 49522 35646 49534 35698
rect 49586 35646 49598 35698
rect 37550 35634 37602 35646
rect 47182 35634 47234 35646
rect 52558 35634 52610 35646
rect 52782 35698 52834 35710
rect 52782 35634 52834 35646
rect 53006 35698 53058 35710
rect 53006 35634 53058 35646
rect 53230 35698 53282 35710
rect 53230 35634 53282 35646
rect 53454 35698 53506 35710
rect 55134 35698 55186 35710
rect 54226 35646 54238 35698
rect 54290 35646 54302 35698
rect 53454 35634 53506 35646
rect 55134 35634 55186 35646
rect 26014 35586 26066 35598
rect 10098 35534 10110 35586
rect 10162 35534 10174 35586
rect 12450 35534 12462 35586
rect 12514 35534 12526 35586
rect 15362 35534 15374 35586
rect 15426 35534 15438 35586
rect 17826 35534 17838 35586
rect 17890 35534 17902 35586
rect 26014 35522 26066 35534
rect 32510 35586 32562 35598
rect 46734 35586 46786 35598
rect 38658 35534 38670 35586
rect 38722 35534 38734 35586
rect 43250 35534 43262 35586
rect 43314 35534 43326 35586
rect 52658 35534 52670 35586
rect 52722 35534 52734 35586
rect 54338 35534 54350 35586
rect 54402 35534 54414 35586
rect 32510 35522 32562 35534
rect 46734 35522 46786 35534
rect 1934 35474 1986 35486
rect 34302 35474 34354 35486
rect 25666 35422 25678 35474
rect 25730 35471 25742 35474
rect 26002 35471 26014 35474
rect 25730 35425 26014 35471
rect 25730 35422 25742 35425
rect 26002 35422 26014 35425
rect 26066 35422 26078 35474
rect 1934 35410 1986 35422
rect 34302 35410 34354 35422
rect 36318 35474 36370 35486
rect 36318 35410 36370 35422
rect 1344 35306 58576 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 58576 35306
rect 1344 35220 58576 35254
rect 5518 35138 5570 35150
rect 33294 35138 33346 35150
rect 20066 35086 20078 35138
rect 20130 35086 20142 35138
rect 31266 35086 31278 35138
rect 31330 35086 31342 35138
rect 5518 35074 5570 35086
rect 33294 35074 33346 35086
rect 34078 35138 34130 35150
rect 34078 35074 34130 35086
rect 44942 35138 44994 35150
rect 48850 35086 48862 35138
rect 48914 35086 48926 35138
rect 44942 35074 44994 35086
rect 12910 35026 12962 35038
rect 12910 34962 12962 34974
rect 18062 35026 18114 35038
rect 20750 35026 20802 35038
rect 18722 34974 18734 35026
rect 18786 34974 18798 35026
rect 18062 34962 18114 34974
rect 20750 34962 20802 34974
rect 22318 35026 22370 35038
rect 22318 34962 22370 34974
rect 25902 35026 25954 35038
rect 28702 35026 28754 35038
rect 33854 35026 33906 35038
rect 40574 35026 40626 35038
rect 27346 34974 27358 35026
rect 27410 34974 27422 35026
rect 30930 34974 30942 35026
rect 30994 34974 31006 35026
rect 38098 34974 38110 35026
rect 38162 34974 38174 35026
rect 25902 34962 25954 34974
rect 28702 34962 28754 34974
rect 33854 34962 33906 34974
rect 40574 34962 40626 34974
rect 50318 35026 50370 35038
rect 50318 34962 50370 34974
rect 8990 34914 9042 34926
rect 8642 34862 8654 34914
rect 8706 34862 8718 34914
rect 8990 34850 9042 34862
rect 13470 34914 13522 34926
rect 19406 34914 19458 34926
rect 24222 34914 24274 34926
rect 14802 34862 14814 34914
rect 14866 34862 14878 34914
rect 19618 34862 19630 34914
rect 19682 34862 19694 34914
rect 21858 34862 21870 34914
rect 21922 34862 21934 34914
rect 22754 34862 22766 34914
rect 22818 34862 22830 34914
rect 13470 34850 13522 34862
rect 19406 34850 19458 34862
rect 24222 34850 24274 34862
rect 24782 34914 24834 34926
rect 24782 34850 24834 34862
rect 26350 34914 26402 34926
rect 29150 34914 29202 34926
rect 30494 34914 30546 34926
rect 39118 34914 39170 34926
rect 44830 34914 44882 34926
rect 27234 34862 27246 34914
rect 27298 34862 27310 34914
rect 30258 34862 30270 34914
rect 30322 34862 30334 34914
rect 31042 34862 31054 34914
rect 31106 34862 31118 34914
rect 32274 34862 32286 34914
rect 32338 34862 32350 34914
rect 37314 34862 37326 34914
rect 37378 34862 37390 34914
rect 38210 34862 38222 34914
rect 38274 34862 38286 34914
rect 43362 34862 43374 34914
rect 43426 34862 43438 34914
rect 26350 34850 26402 34862
rect 29150 34850 29202 34862
rect 30494 34850 30546 34862
rect 39118 34850 39170 34862
rect 44830 34850 44882 34862
rect 46846 34914 46898 34926
rect 48078 34914 48130 34926
rect 49422 34914 49474 34926
rect 47506 34862 47518 34914
rect 47570 34862 47582 34914
rect 48738 34862 48750 34914
rect 48802 34862 48814 34914
rect 49186 34862 49198 34914
rect 49250 34862 49262 34914
rect 46846 34850 46898 34862
rect 48078 34850 48130 34862
rect 49422 34850 49474 34862
rect 49758 34914 49810 34926
rect 52658 34862 52670 34914
rect 52722 34862 52734 34914
rect 54674 34862 54686 34914
rect 54738 34862 54750 34914
rect 49758 34850 49810 34862
rect 10446 34802 10498 34814
rect 18398 34802 18450 34814
rect 9426 34750 9438 34802
rect 9490 34750 9502 34802
rect 13794 34750 13806 34802
rect 13858 34750 13870 34802
rect 15026 34750 15038 34802
rect 15090 34750 15102 34802
rect 10446 34738 10498 34750
rect 18398 34738 18450 34750
rect 18622 34802 18674 34814
rect 32734 34802 32786 34814
rect 26674 34750 26686 34802
rect 26738 34750 26750 34802
rect 29474 34750 29486 34802
rect 29538 34750 29550 34802
rect 18622 34738 18674 34750
rect 32734 34738 32786 34750
rect 33518 34802 33570 34814
rect 44942 34802 44994 34814
rect 37202 34750 37214 34802
rect 37266 34750 37278 34802
rect 38546 34750 38558 34802
rect 38610 34750 38622 34802
rect 33518 34738 33570 34750
rect 44942 34738 44994 34750
rect 46510 34802 46562 34814
rect 46510 34738 46562 34750
rect 49870 34802 49922 34814
rect 55806 34802 55858 34814
rect 52770 34750 52782 34802
rect 52834 34750 52846 34802
rect 49870 34738 49922 34750
rect 55806 34738 55858 34750
rect 9774 34690 9826 34702
rect 6290 34638 6302 34690
rect 6354 34638 6366 34690
rect 9774 34626 9826 34638
rect 10110 34690 10162 34702
rect 10110 34626 10162 34638
rect 10894 34690 10946 34702
rect 10894 34626 10946 34638
rect 11342 34690 11394 34702
rect 11342 34626 11394 34638
rect 14254 34690 14306 34702
rect 32846 34690 32898 34702
rect 22978 34638 22990 34690
rect 23042 34638 23054 34690
rect 32050 34638 32062 34690
rect 32114 34638 32126 34690
rect 14254 34626 14306 34638
rect 32846 34626 32898 34638
rect 34190 34690 34242 34702
rect 34190 34626 34242 34638
rect 39454 34690 39506 34702
rect 46622 34690 46674 34702
rect 43586 34638 43598 34690
rect 43650 34638 43662 34690
rect 52882 34638 52894 34690
rect 52946 34638 52958 34690
rect 39454 34626 39506 34638
rect 46622 34626 46674 34638
rect 1344 34522 58576 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 58576 34522
rect 1344 34436 58576 34470
rect 9102 34354 9154 34366
rect 8306 34302 8318 34354
rect 8370 34302 8382 34354
rect 9102 34290 9154 34302
rect 10558 34354 10610 34366
rect 16830 34354 16882 34366
rect 11106 34302 11118 34354
rect 11170 34302 11182 34354
rect 14466 34302 14478 34354
rect 14530 34302 14542 34354
rect 10558 34290 10610 34302
rect 16830 34290 16882 34302
rect 17390 34354 17442 34366
rect 17390 34290 17442 34302
rect 21646 34354 21698 34366
rect 21646 34290 21698 34302
rect 21758 34354 21810 34366
rect 21758 34290 21810 34302
rect 22430 34354 22482 34366
rect 23550 34354 23602 34366
rect 23202 34302 23214 34354
rect 23266 34302 23278 34354
rect 22430 34290 22482 34302
rect 23550 34290 23602 34302
rect 26014 34354 26066 34366
rect 26014 34290 26066 34302
rect 26238 34354 26290 34366
rect 30606 34354 30658 34366
rect 30146 34302 30158 34354
rect 30210 34302 30222 34354
rect 26238 34290 26290 34302
rect 30606 34290 30658 34302
rect 34190 34354 34242 34366
rect 44494 34354 44546 34366
rect 35746 34302 35758 34354
rect 35810 34302 35822 34354
rect 38882 34302 38894 34354
rect 38946 34302 38958 34354
rect 43922 34302 43934 34354
rect 43986 34302 43998 34354
rect 34190 34290 34242 34302
rect 44494 34290 44546 34302
rect 46398 34354 46450 34366
rect 46398 34290 46450 34302
rect 46510 34354 46562 34366
rect 46510 34290 46562 34302
rect 47854 34354 47906 34366
rect 47854 34290 47906 34302
rect 49870 34354 49922 34366
rect 49870 34290 49922 34302
rect 50878 34354 50930 34366
rect 50878 34290 50930 34302
rect 51998 34354 52050 34366
rect 51998 34290 52050 34302
rect 53790 34354 53842 34366
rect 53790 34290 53842 34302
rect 54350 34354 54402 34366
rect 54350 34290 54402 34302
rect 54462 34354 54514 34366
rect 54462 34290 54514 34302
rect 55582 34354 55634 34366
rect 55582 34290 55634 34302
rect 19630 34242 19682 34254
rect 18386 34190 18398 34242
rect 18450 34190 18462 34242
rect 19058 34190 19070 34242
rect 19122 34190 19134 34242
rect 19630 34178 19682 34190
rect 25678 34242 25730 34254
rect 33630 34242 33682 34254
rect 40014 34242 40066 34254
rect 29250 34190 29262 34242
rect 29314 34190 29326 34242
rect 34850 34190 34862 34242
rect 34914 34190 34926 34242
rect 39218 34190 39230 34242
rect 39282 34190 39294 34242
rect 25678 34178 25730 34190
rect 33630 34178 33682 34190
rect 40014 34178 40066 34190
rect 40350 34242 40402 34254
rect 40350 34178 40402 34190
rect 45390 34242 45442 34254
rect 45390 34178 45442 34190
rect 46846 34242 46898 34254
rect 46846 34178 46898 34190
rect 46958 34242 47010 34254
rect 46958 34178 47010 34190
rect 47630 34242 47682 34254
rect 47630 34178 47682 34190
rect 50654 34242 50706 34254
rect 54238 34242 54290 34254
rect 52994 34190 53006 34242
rect 53058 34190 53070 34242
rect 50654 34178 50706 34190
rect 54238 34178 54290 34190
rect 55246 34242 55298 34254
rect 55246 34178 55298 34190
rect 9550 34130 9602 34142
rect 17950 34130 18002 34142
rect 19518 34130 19570 34142
rect 5506 34078 5518 34130
rect 5570 34078 5582 34130
rect 6066 34078 6078 34130
rect 6130 34078 6142 34130
rect 13682 34078 13694 34130
rect 13746 34078 13758 34130
rect 14130 34078 14142 34130
rect 14194 34078 14206 34130
rect 14690 34078 14702 34130
rect 14754 34078 14766 34130
rect 18722 34078 18734 34130
rect 18786 34078 18798 34130
rect 9550 34066 9602 34078
rect 17950 34066 18002 34078
rect 19518 34066 19570 34078
rect 19742 34130 19794 34142
rect 21086 34130 21138 34142
rect 19842 34078 19854 34130
rect 19906 34078 19918 34130
rect 19742 34066 19794 34078
rect 21086 34066 21138 34078
rect 21310 34130 21362 34142
rect 21310 34066 21362 34078
rect 21534 34130 21586 34142
rect 21534 34066 21586 34078
rect 25566 34130 25618 34142
rect 25566 34066 25618 34078
rect 25902 34130 25954 34142
rect 25902 34066 25954 34078
rect 26350 34130 26402 34142
rect 41022 34130 41074 34142
rect 46286 34130 46338 34142
rect 29698 34078 29710 34130
rect 29762 34078 29774 34130
rect 30034 34078 30046 34130
rect 30098 34078 30110 34130
rect 34738 34078 34750 34130
rect 34802 34078 34814 34130
rect 36306 34078 36318 34130
rect 36370 34078 36382 34130
rect 37874 34078 37886 34130
rect 37938 34078 37950 34130
rect 38658 34078 38670 34130
rect 38722 34078 38734 34130
rect 39442 34078 39454 34130
rect 39506 34078 39518 34130
rect 41346 34078 41358 34130
rect 41410 34078 41422 34130
rect 45154 34078 45166 34130
rect 45218 34078 45230 34130
rect 45938 34078 45950 34130
rect 46002 34078 46014 34130
rect 26350 34066 26402 34078
rect 41022 34066 41074 34078
rect 46286 34066 46338 34078
rect 49646 34130 49698 34142
rect 49646 34066 49698 34078
rect 50094 34130 50146 34142
rect 50094 34066 50146 34078
rect 50206 34130 50258 34142
rect 50206 34066 50258 34078
rect 50766 34130 50818 34142
rect 50766 34066 50818 34078
rect 52446 34130 52498 34142
rect 52446 34066 52498 34078
rect 15262 34018 15314 34030
rect 51886 34018 51938 34030
rect 9986 33966 9998 34018
rect 10050 33966 10062 34018
rect 31042 33966 31054 34018
rect 31106 33966 31118 34018
rect 47954 33966 47966 34018
rect 48018 33966 48030 34018
rect 15262 33954 15314 33966
rect 51886 33954 51938 33966
rect 20190 33906 20242 33918
rect 20190 33842 20242 33854
rect 20862 33906 20914 33918
rect 20862 33842 20914 33854
rect 46958 33906 47010 33918
rect 46958 33842 47010 33854
rect 1344 33738 58576 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 58576 33738
rect 1344 33652 58576 33686
rect 14030 33570 14082 33582
rect 14030 33506 14082 33518
rect 19518 33570 19570 33582
rect 19518 33506 19570 33518
rect 24670 33570 24722 33582
rect 24670 33506 24722 33518
rect 25230 33570 25282 33582
rect 25230 33506 25282 33518
rect 26350 33570 26402 33582
rect 26350 33506 26402 33518
rect 26462 33570 26514 33582
rect 26462 33506 26514 33518
rect 37438 33570 37490 33582
rect 37438 33506 37490 33518
rect 49310 33570 49362 33582
rect 49310 33506 49362 33518
rect 51438 33570 51490 33582
rect 51438 33506 51490 33518
rect 8318 33458 8370 33470
rect 8318 33394 8370 33406
rect 18510 33458 18562 33470
rect 18510 33394 18562 33406
rect 19294 33458 19346 33470
rect 19294 33394 19346 33406
rect 21534 33458 21586 33470
rect 21534 33394 21586 33406
rect 22990 33458 23042 33470
rect 22990 33394 23042 33406
rect 23550 33458 23602 33470
rect 23550 33394 23602 33406
rect 27582 33458 27634 33470
rect 49982 33458 50034 33470
rect 45154 33406 45166 33458
rect 45218 33406 45230 33458
rect 27582 33394 27634 33406
rect 49982 33394 50034 33406
rect 50766 33458 50818 33470
rect 57934 33458 57986 33470
rect 52770 33406 52782 33458
rect 52834 33406 52846 33458
rect 50766 33394 50818 33406
rect 57934 33394 57986 33406
rect 12014 33346 12066 33358
rect 17502 33346 17554 33358
rect 11666 33294 11678 33346
rect 11730 33294 11742 33346
rect 17154 33294 17166 33346
rect 17218 33294 17230 33346
rect 12014 33282 12066 33294
rect 17502 33282 17554 33294
rect 18846 33346 18898 33358
rect 18846 33282 18898 33294
rect 19742 33346 19794 33358
rect 19742 33282 19794 33294
rect 20078 33346 20130 33358
rect 20078 33282 20130 33294
rect 21982 33346 22034 33358
rect 21982 33282 22034 33294
rect 22654 33346 22706 33358
rect 22654 33282 22706 33294
rect 24446 33346 24498 33358
rect 24446 33282 24498 33294
rect 25006 33346 25058 33358
rect 25006 33282 25058 33294
rect 25678 33346 25730 33358
rect 25678 33282 25730 33294
rect 25902 33346 25954 33358
rect 25902 33282 25954 33294
rect 26238 33346 26290 33358
rect 26238 33282 26290 33294
rect 26686 33346 26738 33358
rect 40910 33346 40962 33358
rect 43038 33346 43090 33358
rect 47182 33346 47234 33358
rect 36194 33294 36206 33346
rect 36258 33294 36270 33346
rect 40450 33294 40462 33346
rect 40514 33294 40526 33346
rect 42466 33294 42478 33346
rect 42530 33294 42542 33346
rect 43698 33294 43710 33346
rect 43762 33294 43774 33346
rect 45266 33294 45278 33346
rect 45330 33294 45342 33346
rect 46498 33294 46510 33346
rect 46562 33294 46574 33346
rect 26686 33282 26738 33294
rect 40910 33282 40962 33294
rect 43038 33282 43090 33294
rect 47182 33282 47234 33294
rect 47518 33346 47570 33358
rect 47518 33282 47570 33294
rect 48638 33346 48690 33358
rect 48638 33282 48690 33294
rect 49534 33346 49586 33358
rect 52994 33294 53006 33346
rect 53058 33294 53070 33346
rect 55570 33294 55582 33346
rect 55634 33294 55646 33346
rect 49534 33282 49586 33294
rect 1710 33234 1762 33246
rect 1710 33170 1762 33182
rect 2046 33234 2098 33246
rect 2046 33170 2098 33182
rect 8542 33234 8594 33246
rect 22094 33234 22146 33246
rect 20402 33182 20414 33234
rect 20466 33182 20478 33234
rect 8542 33170 8594 33182
rect 22094 33170 22146 33182
rect 27022 33234 27074 33246
rect 43150 33234 43202 33246
rect 36418 33182 36430 33234
rect 36482 33182 36494 33234
rect 27022 33170 27074 33182
rect 43150 33170 43202 33182
rect 48190 33234 48242 33246
rect 48190 33170 48242 33182
rect 48526 33234 48578 33246
rect 48526 33170 48578 33182
rect 49758 33234 49810 33246
rect 49758 33170 49810 33182
rect 50094 33234 50146 33246
rect 50094 33170 50146 33182
rect 50654 33234 50706 33246
rect 50654 33170 50706 33182
rect 50878 33234 50930 33246
rect 50878 33170 50930 33182
rect 51326 33234 51378 33246
rect 51326 33170 51378 33182
rect 53678 33234 53730 33246
rect 53678 33170 53730 33182
rect 54014 33234 54066 33246
rect 54014 33170 54066 33182
rect 54350 33234 54402 33246
rect 54350 33170 54402 33182
rect 2494 33122 2546 33134
rect 12574 33122 12626 33134
rect 9090 33070 9102 33122
rect 9154 33070 9166 33122
rect 2494 33058 2546 33070
rect 12574 33058 12626 33070
rect 13582 33122 13634 33134
rect 18958 33122 19010 33134
rect 14578 33070 14590 33122
rect 14642 33070 14654 33122
rect 13582 33058 13634 33070
rect 18958 33058 19010 33070
rect 19070 33122 19122 33134
rect 19070 33058 19122 33070
rect 22206 33122 22258 33134
rect 22206 33058 22258 33070
rect 23998 33122 24050 33134
rect 23998 33058 24050 33070
rect 24334 33122 24386 33134
rect 24334 33058 24386 33070
rect 26910 33122 26962 33134
rect 26910 33058 26962 33070
rect 28590 33122 28642 33134
rect 28590 33058 28642 33070
rect 29486 33122 29538 33134
rect 30270 33122 30322 33134
rect 29810 33070 29822 33122
rect 29874 33070 29886 33122
rect 29486 33058 29538 33070
rect 30270 33058 30322 33070
rect 34302 33122 34354 33134
rect 43486 33122 43538 33134
rect 37986 33070 37998 33122
rect 38050 33070 38062 33122
rect 34302 33058 34354 33070
rect 43486 33058 43538 33070
rect 47630 33122 47682 33134
rect 47630 33058 47682 33070
rect 47854 33122 47906 33134
rect 47854 33058 47906 33070
rect 48302 33122 48354 33134
rect 48302 33058 48354 33070
rect 48974 33122 49026 33134
rect 48974 33058 49026 33070
rect 49198 33122 49250 33134
rect 49198 33058 49250 33070
rect 51438 33122 51490 33134
rect 51438 33058 51490 33070
rect 1344 32954 58576 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 58576 32954
rect 1344 32868 58576 32902
rect 19630 32786 19682 32798
rect 19630 32722 19682 32734
rect 20526 32786 20578 32798
rect 20526 32722 20578 32734
rect 22766 32786 22818 32798
rect 22766 32722 22818 32734
rect 22990 32786 23042 32798
rect 22990 32722 23042 32734
rect 24782 32786 24834 32798
rect 24782 32722 24834 32734
rect 25454 32786 25506 32798
rect 29822 32786 29874 32798
rect 37214 32786 37266 32798
rect 29250 32734 29262 32786
rect 29314 32734 29326 32786
rect 36642 32734 36654 32786
rect 36706 32734 36718 32786
rect 25454 32722 25506 32734
rect 29822 32722 29874 32734
rect 37214 32722 37266 32734
rect 43150 32786 43202 32798
rect 43150 32722 43202 32734
rect 43710 32786 43762 32798
rect 48078 32786 48130 32798
rect 47506 32734 47518 32786
rect 47570 32734 47582 32786
rect 50306 32734 50318 32786
rect 50370 32734 50382 32786
rect 43710 32722 43762 32734
rect 48078 32722 48130 32734
rect 19854 32674 19906 32686
rect 19854 32610 19906 32622
rect 23438 32674 23490 32686
rect 23438 32610 23490 32622
rect 25230 32674 25282 32686
rect 38110 32674 38162 32686
rect 43598 32674 43650 32686
rect 37762 32622 37774 32674
rect 37826 32622 37838 32674
rect 38434 32622 38446 32674
rect 38498 32622 38510 32674
rect 25230 32610 25282 32622
rect 38110 32610 38162 32622
rect 43598 32610 43650 32622
rect 43934 32674 43986 32686
rect 43934 32610 43986 32622
rect 46958 32674 47010 32686
rect 46958 32610 47010 32622
rect 47966 32674 48018 32686
rect 47966 32610 48018 32622
rect 49646 32674 49698 32686
rect 49646 32610 49698 32622
rect 19966 32562 20018 32574
rect 16706 32510 16718 32562
rect 16770 32510 16782 32562
rect 19966 32498 20018 32510
rect 22654 32562 22706 32574
rect 22654 32498 22706 32510
rect 23102 32562 23154 32574
rect 23102 32498 23154 32510
rect 25790 32562 25842 32574
rect 25790 32498 25842 32510
rect 26126 32562 26178 32574
rect 47182 32562 47234 32574
rect 26674 32510 26686 32562
rect 26738 32510 26750 32562
rect 30146 32510 30158 32562
rect 30210 32510 30222 32562
rect 33618 32510 33630 32562
rect 33682 32510 33694 32562
rect 34066 32510 34078 32562
rect 34130 32510 34142 32562
rect 37538 32510 37550 32562
rect 37602 32510 37614 32562
rect 26126 32498 26178 32510
rect 47182 32498 47234 32510
rect 48302 32562 48354 32574
rect 48302 32498 48354 32510
rect 49758 32562 49810 32574
rect 49758 32498 49810 32510
rect 49870 32562 49922 32574
rect 49870 32498 49922 32510
rect 1822 32450 1874 32462
rect 25566 32450 25618 32462
rect 11778 32398 11790 32450
rect 11842 32398 11854 32450
rect 1822 32386 1874 32398
rect 25566 32386 25618 32398
rect 30606 32450 30658 32462
rect 30606 32386 30658 32398
rect 23550 32338 23602 32350
rect 23550 32274 23602 32286
rect 1344 32170 58576 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 58576 32170
rect 1344 32084 58576 32118
rect 48862 32002 48914 32014
rect 48862 31938 48914 31950
rect 49198 32002 49250 32014
rect 49198 31938 49250 31950
rect 37102 31890 37154 31902
rect 39342 31890 39394 31902
rect 38994 31838 39006 31890
rect 39058 31838 39070 31890
rect 37102 31826 37154 31838
rect 39342 31826 39394 31838
rect 46174 31890 46226 31902
rect 46174 31826 46226 31838
rect 48638 31890 48690 31902
rect 48638 31826 48690 31838
rect 30046 31778 30098 31790
rect 33742 31778 33794 31790
rect 1810 31726 1822 31778
rect 1874 31726 1886 31778
rect 24434 31726 24446 31778
rect 24498 31726 24510 31778
rect 24994 31726 25006 31778
rect 25058 31726 25070 31778
rect 30482 31726 30494 31778
rect 30546 31726 30558 31778
rect 30046 31714 30098 31726
rect 33742 31714 33794 31726
rect 34190 31778 34242 31790
rect 34190 31714 34242 31726
rect 34302 31778 34354 31790
rect 38658 31726 38670 31778
rect 38722 31726 38734 31778
rect 34302 31714 34354 31726
rect 2382 31666 2434 31678
rect 21310 31666 21362 31678
rect 18498 31614 18510 31666
rect 18562 31614 18574 31666
rect 19282 31614 19294 31666
rect 19346 31614 19358 31666
rect 2382 31602 2434 31614
rect 21310 31602 21362 31614
rect 32734 31666 32786 31678
rect 32734 31602 32786 31614
rect 2046 31554 2098 31566
rect 2046 31490 2098 31502
rect 4622 31554 4674 31566
rect 4622 31490 4674 31502
rect 18174 31554 18226 31566
rect 18174 31490 18226 31502
rect 18958 31554 19010 31566
rect 25902 31554 25954 31566
rect 21970 31502 21982 31554
rect 22034 31502 22046 31554
rect 18958 31490 19010 31502
rect 25902 31490 25954 31502
rect 33518 31554 33570 31566
rect 33518 31490 33570 31502
rect 34078 31554 34130 31566
rect 34078 31490 34130 31502
rect 1344 31386 58576 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 58576 31386
rect 1344 31300 58576 31334
rect 8766 31218 8818 31230
rect 16606 31218 16658 31230
rect 7858 31166 7870 31218
rect 7922 31166 7934 31218
rect 13010 31166 13022 31218
rect 13074 31166 13086 31218
rect 8766 31154 8818 31166
rect 16606 31154 16658 31166
rect 17502 31218 17554 31230
rect 33742 31218 33794 31230
rect 25778 31166 25790 31218
rect 25842 31166 25854 31218
rect 17502 31154 17554 31166
rect 33742 31154 33794 31166
rect 38558 31218 38610 31230
rect 38558 31154 38610 31166
rect 38782 31218 38834 31230
rect 38782 31154 38834 31166
rect 39006 31218 39058 31230
rect 39006 31154 39058 31166
rect 39678 31218 39730 31230
rect 39678 31154 39730 31166
rect 41694 31218 41746 31230
rect 41694 31154 41746 31166
rect 41918 31218 41970 31230
rect 46174 31218 46226 31230
rect 45378 31166 45390 31218
rect 45442 31166 45454 31218
rect 41918 31154 41970 31166
rect 46174 31154 46226 31166
rect 9886 31106 9938 31118
rect 40910 31106 40962 31118
rect 17826 31054 17838 31106
rect 17890 31054 17902 31106
rect 21858 31054 21870 31106
rect 21922 31054 21934 31106
rect 31826 31054 31838 31106
rect 31890 31054 31902 31106
rect 9886 31042 9938 31054
rect 40910 31042 40962 31054
rect 41246 31106 41298 31118
rect 41246 31042 41298 31054
rect 47294 31106 47346 31118
rect 57810 31054 57822 31106
rect 57874 31054 57886 31106
rect 47294 31042 47346 31054
rect 16158 30994 16210 31006
rect 4274 30942 4286 30994
rect 4338 30942 4350 30994
rect 4834 30942 4846 30994
rect 4898 30942 4910 30994
rect 5394 30942 5406 30994
rect 5458 30942 5470 30994
rect 9650 30942 9662 30994
rect 9714 30942 9726 30994
rect 15474 30942 15486 30994
rect 15538 30942 15550 30994
rect 16158 30930 16210 30942
rect 18958 30994 19010 31006
rect 33854 30994 33906 31006
rect 19394 30942 19406 30994
rect 19458 30942 19470 30994
rect 25554 30942 25566 30994
rect 25618 30942 25630 30994
rect 26898 30942 26910 30994
rect 26962 30942 26974 30994
rect 33506 30942 33518 30994
rect 33570 30942 33582 30994
rect 18958 30930 19010 30942
rect 33854 30930 33906 30942
rect 41358 30994 41410 31006
rect 41358 30930 41410 30942
rect 42030 30994 42082 31006
rect 42030 30930 42082 30942
rect 42702 30994 42754 31006
rect 46510 30994 46562 31006
rect 58158 30994 58210 31006
rect 43026 30942 43038 30994
rect 43090 30942 43102 30994
rect 46722 30942 46734 30994
rect 46786 30942 46798 30994
rect 42702 30930 42754 30942
rect 46510 30930 46562 30942
rect 58158 30930 58210 30942
rect 18622 30882 18674 30894
rect 18622 30818 18674 30830
rect 26238 30882 26290 30894
rect 26238 30818 26290 30830
rect 38670 30882 38722 30894
rect 41022 30882 41074 30894
rect 39778 30830 39790 30882
rect 39842 30830 39854 30882
rect 38670 30818 38722 30830
rect 41022 30818 41074 30830
rect 57598 30882 57650 30894
rect 57598 30818 57650 30830
rect 1934 30770 1986 30782
rect 1934 30706 1986 30718
rect 8430 30770 8482 30782
rect 8430 30706 8482 30718
rect 12462 30770 12514 30782
rect 12462 30706 12514 30718
rect 39454 30770 39506 30782
rect 39454 30706 39506 30718
rect 1344 30602 58576 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 58576 30602
rect 1344 30516 58576 30550
rect 38894 30434 38946 30446
rect 38894 30370 38946 30382
rect 42142 30434 42194 30446
rect 42142 30370 42194 30382
rect 23998 30322 24050 30334
rect 21746 30270 21758 30322
rect 21810 30270 21822 30322
rect 23998 30258 24050 30270
rect 32062 30322 32114 30334
rect 32062 30258 32114 30270
rect 11230 30210 11282 30222
rect 4162 30158 4174 30210
rect 4226 30158 4238 30210
rect 10770 30158 10782 30210
rect 10834 30158 10846 30210
rect 11230 30146 11282 30158
rect 11790 30210 11842 30222
rect 17838 30210 17890 30222
rect 13682 30158 13694 30210
rect 13746 30158 13758 30210
rect 17602 30158 17614 30210
rect 17666 30158 17678 30210
rect 11790 30146 11842 30158
rect 17838 30146 17890 30158
rect 19182 30210 19234 30222
rect 19182 30146 19234 30158
rect 19406 30210 19458 30222
rect 23774 30210 23826 30222
rect 19618 30158 19630 30210
rect 19682 30158 19694 30210
rect 20066 30158 20078 30210
rect 20130 30158 20142 30210
rect 21970 30158 21982 30210
rect 22034 30158 22046 30210
rect 19406 30146 19458 30158
rect 23774 30146 23826 30158
rect 24222 30210 24274 30222
rect 24222 30146 24274 30158
rect 25006 30210 25058 30222
rect 33966 30210 34018 30222
rect 45950 30210 46002 30222
rect 25330 30158 25342 30210
rect 25394 30158 25406 30210
rect 32722 30158 32734 30210
rect 32786 30158 32798 30210
rect 38546 30158 38558 30210
rect 38610 30158 38622 30210
rect 25006 30146 25058 30158
rect 33966 30146 34018 30158
rect 45950 30146 46002 30158
rect 5630 30098 5682 30110
rect 2482 30046 2494 30098
rect 2546 30046 2558 30098
rect 5630 30034 5682 30046
rect 5966 30098 6018 30110
rect 5966 30034 6018 30046
rect 8542 30098 8594 30110
rect 8542 30034 8594 30046
rect 13918 30098 13970 30110
rect 13918 30034 13970 30046
rect 16942 30098 16994 30110
rect 16942 30034 16994 30046
rect 18398 30098 18450 30110
rect 18398 30034 18450 30046
rect 18510 30098 18562 30110
rect 18510 30034 18562 30046
rect 21310 30098 21362 30110
rect 21310 30034 21362 30046
rect 30718 30098 30770 30110
rect 30718 30034 30770 30046
rect 31054 30098 31106 30110
rect 31054 30034 31106 30046
rect 31726 30098 31778 30110
rect 33294 30098 33346 30110
rect 44158 30098 44210 30110
rect 32834 30046 32846 30098
rect 32898 30046 32910 30098
rect 40226 30046 40238 30098
rect 40290 30046 40302 30098
rect 31726 30034 31778 30046
rect 33294 30034 33346 30046
rect 44158 30034 44210 30046
rect 44270 30098 44322 30110
rect 44270 30034 44322 30046
rect 45614 30098 45666 30110
rect 45614 30034 45666 30046
rect 45838 30098 45890 30110
rect 45838 30034 45890 30046
rect 7758 29986 7810 29998
rect 7758 29922 7810 29934
rect 18174 29986 18226 29998
rect 18174 29922 18226 29934
rect 21534 29986 21586 29998
rect 21534 29922 21586 29934
rect 21758 29986 21810 29998
rect 21758 29922 21810 29934
rect 22542 29986 22594 29998
rect 22542 29922 22594 29934
rect 24334 29986 24386 29998
rect 24334 29922 24386 29934
rect 24446 29986 24498 29998
rect 28478 29986 28530 29998
rect 27906 29934 27918 29986
rect 27970 29934 27982 29986
rect 24446 29922 24498 29934
rect 28478 29922 28530 29934
rect 33406 29986 33458 29998
rect 33406 29922 33458 29934
rect 33630 29986 33682 29998
rect 33630 29922 33682 29934
rect 37326 29986 37378 29998
rect 39230 29986 39282 29998
rect 43934 29986 43986 29998
rect 37650 29934 37662 29986
rect 37714 29934 37726 29986
rect 39554 29934 39566 29986
rect 39618 29934 39630 29986
rect 37326 29922 37378 29934
rect 39230 29922 39282 29934
rect 43934 29922 43986 29934
rect 1344 29818 58576 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 58576 29818
rect 1344 29732 58576 29766
rect 13694 29650 13746 29662
rect 13694 29586 13746 29598
rect 19070 29650 19122 29662
rect 19070 29586 19122 29598
rect 19966 29650 20018 29662
rect 19966 29586 20018 29598
rect 21982 29650 22034 29662
rect 21982 29586 22034 29598
rect 24670 29650 24722 29662
rect 24670 29586 24722 29598
rect 25342 29650 25394 29662
rect 31614 29650 31666 29662
rect 30818 29598 30830 29650
rect 30882 29598 30894 29650
rect 25342 29586 25394 29598
rect 31614 29586 31666 29598
rect 31726 29650 31778 29662
rect 38446 29650 38498 29662
rect 36306 29598 36318 29650
rect 36370 29598 36382 29650
rect 31726 29586 31778 29598
rect 38446 29586 38498 29598
rect 46398 29650 46450 29662
rect 46398 29586 46450 29598
rect 10110 29538 10162 29550
rect 17950 29538 18002 29550
rect 14018 29486 14030 29538
rect 14082 29486 14094 29538
rect 10110 29474 10162 29486
rect 17950 29474 18002 29486
rect 19854 29538 19906 29550
rect 19854 29474 19906 29486
rect 22206 29538 22258 29550
rect 22206 29474 22258 29486
rect 22318 29538 22370 29550
rect 22318 29474 22370 29486
rect 25230 29538 25282 29550
rect 25230 29474 25282 29486
rect 26238 29538 26290 29550
rect 26238 29474 26290 29486
rect 31950 29538 32002 29550
rect 31950 29474 32002 29486
rect 32062 29538 32114 29550
rect 32062 29474 32114 29486
rect 38334 29538 38386 29550
rect 38334 29474 38386 29486
rect 38782 29538 38834 29550
rect 38782 29474 38834 29486
rect 45614 29538 45666 29550
rect 45614 29474 45666 29486
rect 11006 29426 11058 29438
rect 4274 29374 4286 29426
rect 4338 29374 4350 29426
rect 10546 29374 10558 29426
rect 10610 29374 10622 29426
rect 11006 29362 11058 29374
rect 14366 29426 14418 29438
rect 14366 29362 14418 29374
rect 15598 29426 15650 29438
rect 15598 29362 15650 29374
rect 17614 29426 17666 29438
rect 17614 29362 17666 29374
rect 17838 29426 17890 29438
rect 17838 29362 17890 29374
rect 18174 29426 18226 29438
rect 18174 29362 18226 29374
rect 18398 29426 18450 29438
rect 18398 29362 18450 29374
rect 18846 29426 18898 29438
rect 21646 29426 21698 29438
rect 21186 29374 21198 29426
rect 21250 29374 21262 29426
rect 18846 29362 18898 29374
rect 21646 29362 21698 29374
rect 25454 29426 25506 29438
rect 25454 29362 25506 29374
rect 25678 29426 25730 29438
rect 25678 29362 25730 29374
rect 28142 29426 28194 29438
rect 33182 29426 33234 29438
rect 39118 29426 39170 29438
rect 42702 29426 42754 29438
rect 28578 29374 28590 29426
rect 28642 29374 28654 29426
rect 33730 29374 33742 29426
rect 33794 29374 33806 29426
rect 39442 29374 39454 29426
rect 39506 29374 39518 29426
rect 43250 29374 43262 29426
rect 43314 29374 43326 29426
rect 28142 29362 28194 29374
rect 33182 29362 33234 29374
rect 39118 29362 39170 29374
rect 42702 29362 42754 29374
rect 9774 29314 9826 29326
rect 9774 29250 9826 29262
rect 14926 29314 14978 29326
rect 16718 29314 16770 29326
rect 16034 29262 16046 29314
rect 16098 29262 16110 29314
rect 14926 29250 14978 29262
rect 16718 29250 16770 29262
rect 18622 29314 18674 29326
rect 18622 29250 18674 29262
rect 18958 29314 19010 29326
rect 18958 29250 19010 29262
rect 19742 29314 19794 29326
rect 22878 29314 22930 29326
rect 20738 29262 20750 29314
rect 20802 29262 20814 29314
rect 19742 29250 19794 29262
rect 22878 29250 22930 29262
rect 24222 29314 24274 29326
rect 24222 29250 24274 29262
rect 37886 29314 37938 29326
rect 37886 29250 37938 29262
rect 40238 29314 40290 29326
rect 40238 29250 40290 29262
rect 1934 29202 1986 29214
rect 1934 29138 1986 29150
rect 22318 29202 22370 29214
rect 36878 29202 36930 29214
rect 24210 29150 24222 29202
rect 24274 29199 24286 29202
rect 24434 29199 24446 29202
rect 24274 29153 24446 29199
rect 24274 29150 24286 29153
rect 24434 29150 24446 29153
rect 24498 29199 24510 29202
rect 24770 29199 24782 29202
rect 24498 29153 24782 29199
rect 24498 29150 24510 29153
rect 24770 29150 24782 29153
rect 24834 29150 24846 29202
rect 22318 29138 22370 29150
rect 36878 29138 36930 29150
rect 39790 29202 39842 29214
rect 39790 29138 39842 29150
rect 1344 29034 58576 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 58576 29034
rect 1344 28948 58576 28982
rect 31390 28866 31442 28878
rect 31390 28802 31442 28814
rect 1934 28754 1986 28766
rect 18622 28754 18674 28766
rect 15026 28702 15038 28754
rect 15090 28702 15102 28754
rect 1934 28690 1986 28702
rect 18622 28690 18674 28702
rect 19294 28754 19346 28766
rect 19294 28690 19346 28702
rect 21422 28754 21474 28766
rect 21422 28690 21474 28702
rect 24222 28754 24274 28766
rect 33070 28754 33122 28766
rect 25218 28702 25230 28754
rect 25282 28702 25294 28754
rect 24222 28690 24274 28702
rect 33070 28690 33122 28702
rect 33966 28754 34018 28766
rect 33966 28690 34018 28702
rect 6974 28642 7026 28654
rect 4274 28590 4286 28642
rect 4338 28590 4350 28642
rect 6974 28578 7026 28590
rect 9774 28642 9826 28654
rect 9774 28578 9826 28590
rect 10110 28642 10162 28654
rect 13470 28642 13522 28654
rect 10546 28590 10558 28642
rect 10610 28590 10622 28642
rect 12002 28590 12014 28642
rect 12066 28590 12078 28642
rect 10110 28578 10162 28590
rect 13470 28578 13522 28590
rect 13582 28642 13634 28654
rect 13582 28578 13634 28590
rect 13918 28642 13970 28654
rect 15486 28642 15538 28654
rect 14690 28590 14702 28642
rect 14754 28590 14766 28642
rect 13918 28578 13970 28590
rect 15486 28578 15538 28590
rect 16382 28642 16434 28654
rect 16382 28578 16434 28590
rect 17838 28642 17890 28654
rect 17838 28578 17890 28590
rect 19742 28642 19794 28654
rect 19742 28578 19794 28590
rect 21310 28642 21362 28654
rect 21310 28578 21362 28590
rect 21982 28642 22034 28654
rect 21982 28578 22034 28590
rect 22318 28642 22370 28654
rect 22318 28578 22370 28590
rect 22766 28642 22818 28654
rect 25566 28642 25618 28654
rect 24546 28590 24558 28642
rect 24610 28590 24622 28642
rect 22766 28578 22818 28590
rect 25566 28578 25618 28590
rect 26126 28642 26178 28654
rect 26126 28578 26178 28590
rect 29486 28642 29538 28654
rect 29486 28578 29538 28590
rect 31054 28642 31106 28654
rect 37214 28642 37266 28654
rect 31826 28590 31838 28642
rect 31890 28590 31902 28642
rect 33506 28590 33518 28642
rect 33570 28590 33582 28642
rect 31054 28578 31106 28590
rect 37214 28578 37266 28590
rect 37326 28642 37378 28654
rect 37326 28578 37378 28590
rect 37774 28642 37826 28654
rect 37774 28578 37826 28590
rect 38222 28642 38274 28654
rect 38222 28578 38274 28590
rect 11566 28530 11618 28542
rect 11566 28466 11618 28478
rect 16046 28530 16098 28542
rect 20526 28530 20578 28542
rect 16706 28478 16718 28530
rect 16770 28478 16782 28530
rect 18162 28478 18174 28530
rect 18226 28478 18238 28530
rect 16046 28466 16098 28478
rect 20526 28466 20578 28478
rect 20638 28530 20690 28542
rect 29150 28530 29202 28542
rect 33182 28530 33234 28542
rect 24658 28478 24670 28530
rect 24722 28478 24734 28530
rect 32162 28478 32174 28530
rect 32226 28478 32238 28530
rect 20638 28466 20690 28478
rect 29150 28466 29202 28478
rect 33182 28466 33234 28478
rect 37102 28530 37154 28542
rect 37102 28466 37154 28478
rect 38558 28530 38610 28542
rect 38558 28466 38610 28478
rect 9214 28418 9266 28430
rect 7298 28366 7310 28418
rect 7362 28366 7374 28418
rect 9214 28354 9266 28366
rect 13022 28418 13074 28430
rect 17614 28418 17666 28430
rect 14242 28366 14254 28418
rect 14306 28366 14318 28418
rect 13022 28354 13074 28366
rect 17614 28354 17666 28366
rect 20302 28418 20354 28430
rect 20302 28354 20354 28366
rect 20862 28418 20914 28430
rect 20862 28354 20914 28366
rect 21534 28418 21586 28430
rect 21534 28354 21586 28366
rect 28478 28418 28530 28430
rect 28478 28354 28530 28366
rect 32958 28418 33010 28430
rect 32958 28354 33010 28366
rect 58158 28418 58210 28430
rect 58158 28354 58210 28366
rect 1344 28250 58576 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 58576 28250
rect 1344 28164 58576 28198
rect 8878 28082 8930 28094
rect 7298 28030 7310 28082
rect 7362 28030 7374 28082
rect 8878 28018 8930 28030
rect 15598 28082 15650 28094
rect 15598 28018 15650 28030
rect 18958 28082 19010 28094
rect 18958 28018 19010 28030
rect 24670 28082 24722 28094
rect 24670 28018 24722 28030
rect 26910 28082 26962 28094
rect 26910 28018 26962 28030
rect 27694 28082 27746 28094
rect 27694 28018 27746 28030
rect 29038 28082 29090 28094
rect 29038 28018 29090 28030
rect 29822 28082 29874 28094
rect 29822 28018 29874 28030
rect 30830 28082 30882 28094
rect 30830 28018 30882 28030
rect 32622 28082 32674 28094
rect 32622 28018 32674 28030
rect 35534 28082 35586 28094
rect 43922 28030 43934 28082
rect 43986 28030 43998 28082
rect 35534 28018 35586 28030
rect 8430 27970 8482 27982
rect 8430 27906 8482 27918
rect 9550 27970 9602 27982
rect 9550 27906 9602 27918
rect 9886 27970 9938 27982
rect 16270 27970 16322 27982
rect 13234 27918 13246 27970
rect 13298 27918 13310 27970
rect 13794 27918 13806 27970
rect 13858 27918 13870 27970
rect 9886 27906 9938 27918
rect 16270 27906 16322 27918
rect 26126 27970 26178 27982
rect 26126 27906 26178 27918
rect 35646 27970 35698 27982
rect 38222 27970 38274 27982
rect 36418 27918 36430 27970
rect 36482 27918 36494 27970
rect 35646 27906 35698 27918
rect 38222 27906 38274 27918
rect 38558 27970 38610 27982
rect 38558 27906 38610 27918
rect 38670 27970 38722 27982
rect 38670 27906 38722 27918
rect 4622 27858 4674 27870
rect 10558 27858 10610 27870
rect 5058 27806 5070 27858
rect 5122 27806 5134 27858
rect 4622 27794 4674 27806
rect 10558 27794 10610 27806
rect 10782 27858 10834 27870
rect 10782 27794 10834 27806
rect 11006 27858 11058 27870
rect 11006 27794 11058 27806
rect 11230 27858 11282 27870
rect 11230 27794 11282 27806
rect 12350 27858 12402 27870
rect 12350 27794 12402 27806
rect 17390 27858 17442 27870
rect 28030 27858 28082 27870
rect 23538 27806 23550 27858
rect 23602 27806 23614 27858
rect 25666 27806 25678 27858
rect 25730 27806 25742 27858
rect 17390 27794 17442 27806
rect 28030 27794 28082 27806
rect 40798 27858 40850 27870
rect 41346 27806 41358 27858
rect 41410 27806 41422 27858
rect 40798 27794 40850 27806
rect 12126 27746 12178 27758
rect 12126 27682 12178 27694
rect 14366 27746 14418 27758
rect 16830 27746 16882 27758
rect 15138 27694 15150 27746
rect 15202 27694 15214 27746
rect 14366 27682 14418 27694
rect 16830 27682 16882 27694
rect 17950 27746 18002 27758
rect 19518 27746 19570 27758
rect 18498 27694 18510 27746
rect 18562 27694 18574 27746
rect 17950 27682 18002 27694
rect 19518 27682 19570 27694
rect 19854 27746 19906 27758
rect 19854 27682 19906 27694
rect 23998 27746 24050 27758
rect 25330 27694 25342 27746
rect 25394 27694 25406 27746
rect 26450 27694 26462 27746
rect 26514 27694 26526 27746
rect 28466 27694 28478 27746
rect 28530 27694 28542 27746
rect 23998 27682 24050 27694
rect 8094 27634 8146 27646
rect 8094 27570 8146 27582
rect 8318 27634 8370 27646
rect 8318 27570 8370 27582
rect 11678 27634 11730 27646
rect 14030 27634 14082 27646
rect 12674 27582 12686 27634
rect 12738 27582 12750 27634
rect 11678 27570 11730 27582
rect 14030 27570 14082 27582
rect 35534 27634 35586 27646
rect 35534 27570 35586 27582
rect 38558 27634 38610 27646
rect 38558 27570 38610 27582
rect 44494 27634 44546 27646
rect 44494 27570 44546 27582
rect 1344 27466 58576 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 58576 27466
rect 1344 27380 58576 27414
rect 1934 27298 1986 27310
rect 16270 27298 16322 27310
rect 11218 27246 11230 27298
rect 11282 27246 11294 27298
rect 14242 27246 14254 27298
rect 14306 27246 14318 27298
rect 1934 27234 1986 27246
rect 9550 27186 9602 27198
rect 7634 27134 7646 27186
rect 7698 27134 7710 27186
rect 8530 27134 8542 27186
rect 8594 27134 8606 27186
rect 14018 27134 14030 27186
rect 14082 27183 14094 27186
rect 14257 27183 14303 27246
rect 16270 27234 16322 27246
rect 27694 27298 27746 27310
rect 27694 27234 27746 27246
rect 14082 27137 14303 27183
rect 16606 27186 16658 27198
rect 14082 27134 14094 27137
rect 9550 27122 9602 27134
rect 16606 27122 16658 27134
rect 19854 27186 19906 27198
rect 22318 27186 22370 27198
rect 21746 27134 21758 27186
rect 21810 27134 21822 27186
rect 19854 27122 19906 27134
rect 22318 27122 22370 27134
rect 22766 27186 22818 27198
rect 27582 27186 27634 27198
rect 35758 27186 35810 27198
rect 24210 27134 24222 27186
rect 24274 27134 24286 27186
rect 28466 27134 28478 27186
rect 28530 27134 28542 27186
rect 29362 27134 29374 27186
rect 29426 27134 29438 27186
rect 22766 27122 22818 27134
rect 27582 27122 27634 27134
rect 35758 27122 35810 27134
rect 37102 27186 37154 27198
rect 42578 27134 42590 27186
rect 42642 27134 42654 27186
rect 37102 27122 37154 27134
rect 10670 27074 10722 27086
rect 4274 27022 4286 27074
rect 4338 27022 4350 27074
rect 6626 27022 6638 27074
rect 6690 27022 6702 27074
rect 7298 27022 7310 27074
rect 7362 27022 7374 27074
rect 8194 27022 8206 27074
rect 8258 27022 8270 27074
rect 10434 27022 10446 27074
rect 10498 27022 10510 27074
rect 10670 27010 10722 27022
rect 10782 27074 10834 27086
rect 10782 27010 10834 27022
rect 11566 27074 11618 27086
rect 11566 27010 11618 27022
rect 12910 27074 12962 27086
rect 14478 27074 14530 27086
rect 15710 27074 15762 27086
rect 14018 27022 14030 27074
rect 14082 27022 14094 27074
rect 14914 27022 14926 27074
rect 14978 27022 14990 27074
rect 12910 27010 12962 27022
rect 14478 27010 14530 27022
rect 15710 27010 15762 27022
rect 17166 27074 17218 27086
rect 18062 27074 18114 27086
rect 28030 27074 28082 27086
rect 30158 27074 30210 27086
rect 17602 27022 17614 27074
rect 17666 27022 17678 27074
rect 18386 27022 18398 27074
rect 18450 27022 18462 27074
rect 23202 27022 23214 27074
rect 23266 27022 23278 27074
rect 25442 27022 25454 27074
rect 25506 27022 25518 27074
rect 27234 27022 27246 27074
rect 27298 27022 27310 27074
rect 29138 27022 29150 27074
rect 29202 27022 29214 27074
rect 17166 27010 17218 27022
rect 18062 27010 18114 27022
rect 28030 27010 28082 27022
rect 30158 27010 30210 27022
rect 31278 27074 31330 27086
rect 36990 27074 37042 27086
rect 31714 27022 31726 27074
rect 31778 27022 31790 27074
rect 35186 27022 35198 27074
rect 35250 27022 35262 27074
rect 31278 27010 31330 27022
rect 36990 27010 37042 27022
rect 38782 27074 38834 27086
rect 43038 27074 43090 27086
rect 39218 27022 39230 27074
rect 39282 27022 39294 27074
rect 38782 27010 38834 27022
rect 43038 27010 43090 27022
rect 43486 27074 43538 27086
rect 43486 27010 43538 27022
rect 8990 26962 9042 26974
rect 8990 26898 9042 26910
rect 12126 26962 12178 26974
rect 12126 26898 12178 26910
rect 13470 26962 13522 26974
rect 13470 26898 13522 26910
rect 13582 26962 13634 26974
rect 13582 26898 13634 26910
rect 13694 26962 13746 26974
rect 13694 26898 13746 26910
rect 16046 26962 16098 26974
rect 16046 26898 16098 26910
rect 18846 26962 18898 26974
rect 18846 26898 18898 26910
rect 20414 26962 20466 26974
rect 20414 26898 20466 26910
rect 21310 26962 21362 26974
rect 30718 26962 30770 26974
rect 23538 26910 23550 26962
rect 23602 26910 23614 26962
rect 25778 26910 25790 26962
rect 25842 26910 25854 26962
rect 27122 26910 27134 26962
rect 27186 26910 27198 26962
rect 29250 26910 29262 26962
rect 29314 26910 29326 26962
rect 21310 26898 21362 26910
rect 30718 26898 30770 26910
rect 33966 26962 34018 26974
rect 37438 26962 37490 26974
rect 34962 26910 34974 26962
rect 35026 26910 35038 26962
rect 33966 26898 34018 26910
rect 37438 26898 37490 26910
rect 41470 26962 41522 26974
rect 41470 26898 41522 26910
rect 6862 26850 6914 26862
rect 6862 26786 6914 26798
rect 19406 26850 19458 26862
rect 19406 26786 19458 26798
rect 20750 26850 20802 26862
rect 20750 26786 20802 26798
rect 34750 26850 34802 26862
rect 34750 26786 34802 26798
rect 37214 26850 37266 26862
rect 37214 26786 37266 26798
rect 42254 26850 42306 26862
rect 42254 26786 42306 26798
rect 58158 26850 58210 26862
rect 58158 26786 58210 26798
rect 1344 26682 58576 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 58576 26682
rect 1344 26596 58576 26630
rect 1710 26514 1762 26526
rect 39790 26514 39842 26526
rect 16258 26462 16270 26514
rect 16322 26462 16334 26514
rect 45154 26462 45166 26514
rect 45218 26462 45230 26514
rect 1710 26450 1762 26462
rect 39790 26450 39842 26462
rect 20526 26402 20578 26414
rect 39230 26402 39282 26414
rect 5058 26350 5070 26402
rect 5122 26350 5134 26402
rect 6066 26350 6078 26402
rect 6130 26350 6142 26402
rect 15586 26350 15598 26402
rect 15650 26350 15662 26402
rect 24322 26350 24334 26402
rect 24386 26350 24398 26402
rect 27682 26350 27694 26402
rect 27746 26350 27758 26402
rect 20526 26338 20578 26350
rect 39230 26338 39282 26350
rect 58158 26402 58210 26414
rect 58158 26338 58210 26350
rect 8094 26290 8146 26302
rect 4834 26238 4846 26290
rect 4898 26238 4910 26290
rect 8094 26226 8146 26238
rect 10110 26290 10162 26302
rect 14254 26290 14306 26302
rect 18286 26290 18338 26302
rect 10322 26238 10334 26290
rect 10386 26238 10398 26290
rect 12226 26238 12238 26290
rect 12290 26238 12302 26290
rect 13794 26238 13806 26290
rect 13858 26238 13870 26290
rect 14690 26238 14702 26290
rect 14754 26238 14766 26290
rect 15250 26238 15262 26290
rect 15314 26238 15326 26290
rect 16146 26238 16158 26290
rect 16210 26238 16222 26290
rect 10110 26226 10162 26238
rect 14254 26226 14306 26238
rect 18286 26226 18338 26238
rect 18622 26290 18674 26302
rect 18622 26226 18674 26238
rect 19070 26290 19122 26302
rect 31054 26290 31106 26302
rect 38894 26290 38946 26302
rect 20178 26238 20190 26290
rect 20242 26238 20254 26290
rect 21522 26238 21534 26290
rect 21586 26238 21598 26290
rect 22194 26238 22206 26290
rect 22258 26238 22270 26290
rect 22978 26238 22990 26290
rect 23042 26238 23054 26290
rect 24434 26238 24446 26290
rect 24498 26238 24510 26290
rect 26450 26238 26462 26290
rect 26514 26238 26526 26290
rect 28242 26238 28254 26290
rect 28306 26238 28318 26290
rect 29138 26238 29150 26290
rect 29202 26238 29214 26290
rect 30370 26238 30382 26290
rect 30434 26238 30446 26290
rect 31266 26238 31278 26290
rect 31330 26238 31342 26290
rect 19070 26226 19122 26238
rect 31054 26226 31106 26238
rect 38894 26226 38946 26238
rect 42254 26290 42306 26302
rect 42802 26238 42814 26290
rect 42866 26238 42878 26290
rect 42254 26226 42306 26238
rect 6862 26178 6914 26190
rect 5954 26126 5966 26178
rect 6018 26126 6030 26178
rect 6862 26114 6914 26126
rect 8654 26178 8706 26190
rect 8654 26114 8706 26126
rect 9774 26178 9826 26190
rect 12686 26178 12738 26190
rect 16830 26178 16882 26190
rect 19406 26178 19458 26190
rect 11666 26126 11678 26178
rect 11730 26126 11742 26178
rect 13458 26126 13470 26178
rect 13522 26126 13534 26178
rect 17826 26126 17838 26178
rect 17890 26126 17902 26178
rect 9774 26114 9826 26126
rect 12686 26114 12738 26126
rect 16830 26114 16882 26126
rect 19406 26114 19458 26126
rect 19742 26178 19794 26190
rect 19742 26114 19794 26126
rect 20862 26178 20914 26190
rect 23762 26126 23774 26178
rect 23826 26126 23838 26178
rect 26338 26126 26350 26178
rect 26402 26126 26414 26178
rect 20862 26114 20914 26126
rect 2158 26066 2210 26078
rect 45950 26066 46002 26078
rect 13682 26014 13694 26066
rect 13746 26014 13758 26066
rect 28466 26014 28478 26066
rect 28530 26014 28542 26066
rect 31602 26014 31614 26066
rect 31666 26014 31678 26066
rect 2158 26002 2210 26014
rect 45950 26002 46002 26014
rect 1344 25898 58576 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 58576 25898
rect 1344 25812 58576 25846
rect 7086 25730 7138 25742
rect 7086 25666 7138 25678
rect 7422 25730 7474 25742
rect 7422 25666 7474 25678
rect 9326 25730 9378 25742
rect 42814 25730 42866 25742
rect 11330 25678 11342 25730
rect 11394 25678 11406 25730
rect 30482 25678 30494 25730
rect 30546 25727 30558 25730
rect 31266 25727 31278 25730
rect 30546 25681 31278 25727
rect 30546 25678 30558 25681
rect 31266 25678 31278 25681
rect 31330 25678 31342 25730
rect 9326 25666 9378 25678
rect 42814 25666 42866 25678
rect 11902 25618 11954 25630
rect 17390 25618 17442 25630
rect 15362 25566 15374 25618
rect 15426 25566 15438 25618
rect 16482 25566 16494 25618
rect 16546 25566 16558 25618
rect 11902 25554 11954 25566
rect 17390 25554 17442 25566
rect 21758 25618 21810 25630
rect 30718 25618 30770 25630
rect 22754 25566 22766 25618
rect 22818 25566 22830 25618
rect 25890 25566 25902 25618
rect 25954 25566 25966 25618
rect 28130 25566 28142 25618
rect 28194 25566 28206 25618
rect 21758 25554 21810 25566
rect 30718 25554 30770 25566
rect 31278 25618 31330 25630
rect 31278 25554 31330 25566
rect 31614 25618 31666 25630
rect 31614 25554 31666 25566
rect 32174 25618 32226 25630
rect 32174 25554 32226 25566
rect 36094 25618 36146 25630
rect 36094 25554 36146 25566
rect 42366 25618 42418 25630
rect 42366 25554 42418 25566
rect 57934 25618 57986 25630
rect 57934 25554 57986 25566
rect 5966 25506 6018 25518
rect 5966 25442 6018 25454
rect 9438 25506 9490 25518
rect 10670 25506 10722 25518
rect 12238 25506 12290 25518
rect 9874 25454 9886 25506
rect 9938 25454 9950 25506
rect 10994 25454 11006 25506
rect 11058 25454 11070 25506
rect 9438 25442 9490 25454
rect 10670 25442 10722 25454
rect 12238 25442 12290 25454
rect 12686 25506 12738 25518
rect 12686 25442 12738 25454
rect 13918 25506 13970 25518
rect 22318 25506 22370 25518
rect 14130 25454 14142 25506
rect 14194 25454 14206 25506
rect 15250 25454 15262 25506
rect 15314 25454 15326 25506
rect 15922 25454 15934 25506
rect 15986 25454 15998 25506
rect 17042 25454 17054 25506
rect 17106 25454 17118 25506
rect 17938 25454 17950 25506
rect 18002 25454 18014 25506
rect 20178 25454 20190 25506
rect 20242 25454 20254 25506
rect 13918 25442 13970 25454
rect 22318 25442 22370 25454
rect 23214 25506 23266 25518
rect 23214 25442 23266 25454
rect 23886 25506 23938 25518
rect 31838 25506 31890 25518
rect 25106 25454 25118 25506
rect 25170 25454 25182 25506
rect 26114 25454 26126 25506
rect 26178 25454 26190 25506
rect 28578 25454 28590 25506
rect 28642 25454 28654 25506
rect 29138 25454 29150 25506
rect 29202 25454 29214 25506
rect 30034 25454 30046 25506
rect 30098 25454 30110 25506
rect 23886 25442 23938 25454
rect 31838 25442 31890 25454
rect 34414 25506 34466 25518
rect 38558 25506 38610 25518
rect 35074 25454 35086 25506
rect 35138 25454 35150 25506
rect 35522 25454 35534 25506
rect 35586 25454 35598 25506
rect 37986 25454 37998 25506
rect 38050 25454 38062 25506
rect 34414 25442 34466 25454
rect 38558 25442 38610 25454
rect 43934 25506 43986 25518
rect 46834 25454 46846 25506
rect 46898 25454 46910 25506
rect 55570 25454 55582 25506
rect 55634 25454 55646 25506
rect 43934 25442 43986 25454
rect 6862 25394 6914 25406
rect 5618 25342 5630 25394
rect 5682 25342 5694 25394
rect 6862 25330 6914 25342
rect 9326 25394 9378 25406
rect 9326 25330 9378 25342
rect 10334 25394 10386 25406
rect 10334 25330 10386 25342
rect 12462 25394 12514 25406
rect 12462 25330 12514 25342
rect 12910 25394 12962 25406
rect 12910 25330 12962 25342
rect 13022 25394 13074 25406
rect 17614 25394 17666 25406
rect 15474 25342 15486 25394
rect 15538 25342 15550 25394
rect 16258 25342 16270 25394
rect 16322 25342 16334 25394
rect 13022 25330 13074 25342
rect 17614 25330 17666 25342
rect 17726 25394 17778 25406
rect 21534 25394 21586 25406
rect 35758 25394 35810 25406
rect 38670 25394 38722 25406
rect 19282 25342 19294 25394
rect 19346 25342 19358 25394
rect 29250 25342 29262 25394
rect 29314 25342 29326 25394
rect 37314 25342 37326 25394
rect 37378 25342 37390 25394
rect 17726 25330 17778 25342
rect 21534 25330 21586 25342
rect 35758 25330 35810 25342
rect 38670 25330 38722 25342
rect 42814 25394 42866 25406
rect 42814 25330 42866 25342
rect 42926 25394 42978 25406
rect 42926 25330 42978 25342
rect 43150 25394 43202 25406
rect 43150 25330 43202 25342
rect 43374 25394 43426 25406
rect 43374 25330 43426 25342
rect 43486 25394 43538 25406
rect 47058 25342 47070 25394
rect 47122 25342 47134 25394
rect 43486 25330 43538 25342
rect 8990 25282 9042 25294
rect 8990 25218 9042 25230
rect 13582 25282 13634 25294
rect 13582 25218 13634 25230
rect 18398 25282 18450 25294
rect 18398 25218 18450 25230
rect 18958 25282 19010 25294
rect 36206 25282 36258 25294
rect 24546 25230 24558 25282
rect 24610 25230 24622 25282
rect 30146 25230 30158 25282
rect 30210 25230 30222 25282
rect 34066 25230 34078 25282
rect 34130 25230 34142 25282
rect 18958 25218 19010 25230
rect 36206 25218 36258 25230
rect 36990 25282 37042 25294
rect 36990 25218 37042 25230
rect 1344 25114 58576 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 58576 25114
rect 1344 25028 58576 25062
rect 7422 24946 7474 24958
rect 7422 24882 7474 24894
rect 16158 24946 16210 24958
rect 16158 24882 16210 24894
rect 17502 24946 17554 24958
rect 17502 24882 17554 24894
rect 24670 24946 24722 24958
rect 24670 24882 24722 24894
rect 27470 24946 27522 24958
rect 27470 24882 27522 24894
rect 27806 24946 27858 24958
rect 27806 24882 27858 24894
rect 29262 24946 29314 24958
rect 29262 24882 29314 24894
rect 29710 24946 29762 24958
rect 29710 24882 29762 24894
rect 30606 24946 30658 24958
rect 30606 24882 30658 24894
rect 38894 24946 38946 24958
rect 38894 24882 38946 24894
rect 8990 24834 9042 24846
rect 13022 24834 13074 24846
rect 24110 24834 24162 24846
rect 12002 24782 12014 24834
rect 12066 24782 12078 24834
rect 12674 24782 12686 24834
rect 12738 24782 12750 24834
rect 14914 24782 14926 24834
rect 14978 24782 14990 24834
rect 20962 24782 20974 24834
rect 21026 24782 21038 24834
rect 23426 24782 23438 24834
rect 23490 24782 23502 24834
rect 8990 24770 9042 24782
rect 13022 24770 13074 24782
rect 24110 24770 24162 24782
rect 28366 24834 28418 24846
rect 28366 24770 28418 24782
rect 28702 24834 28754 24846
rect 38782 24834 38834 24846
rect 33394 24782 33406 24834
rect 33458 24782 33470 24834
rect 36082 24782 36094 24834
rect 36146 24782 36158 24834
rect 28702 24770 28754 24782
rect 38782 24770 38834 24782
rect 41358 24834 41410 24846
rect 41358 24770 41410 24782
rect 43262 24834 43314 24846
rect 43262 24770 43314 24782
rect 46846 24834 46898 24846
rect 46846 24770 46898 24782
rect 6078 24722 6130 24734
rect 9550 24722 9602 24734
rect 12910 24722 12962 24734
rect 8530 24670 8542 24722
rect 8594 24670 8606 24722
rect 10098 24670 10110 24722
rect 10162 24670 10174 24722
rect 6078 24658 6130 24670
rect 9550 24658 9602 24670
rect 12910 24658 12962 24670
rect 13470 24722 13522 24734
rect 21870 24722 21922 24734
rect 30942 24722 30994 24734
rect 15810 24670 15822 24722
rect 15874 24670 15886 24722
rect 17826 24670 17838 24722
rect 17890 24670 17902 24722
rect 18386 24670 18398 24722
rect 18450 24670 18462 24722
rect 20178 24670 20190 24722
rect 20242 24670 20254 24722
rect 22418 24670 22430 24722
rect 22482 24670 22494 24722
rect 23202 24670 23214 24722
rect 23266 24670 23278 24722
rect 25554 24670 25566 24722
rect 25618 24670 25630 24722
rect 26562 24670 26574 24722
rect 26626 24670 26638 24722
rect 13470 24658 13522 24670
rect 21870 24658 21922 24670
rect 30942 24658 30994 24670
rect 31166 24722 31218 24734
rect 31166 24658 31218 24670
rect 31838 24722 31890 24734
rect 37886 24722 37938 24734
rect 33170 24670 33182 24722
rect 33234 24670 33246 24722
rect 34962 24670 34974 24722
rect 35026 24670 35038 24722
rect 35522 24670 35534 24722
rect 35586 24670 35598 24722
rect 36866 24670 36878 24722
rect 36930 24670 36942 24722
rect 31838 24658 31890 24670
rect 37886 24658 37938 24670
rect 38110 24722 38162 24734
rect 38110 24658 38162 24670
rect 39118 24722 39170 24734
rect 42242 24670 42254 24722
rect 42306 24670 42318 24722
rect 42690 24670 42702 24722
rect 42754 24670 42766 24722
rect 46162 24670 46174 24722
rect 46226 24670 46238 24722
rect 46610 24670 46622 24722
rect 46674 24670 46686 24722
rect 39118 24658 39170 24670
rect 6638 24610 6690 24622
rect 26910 24610 26962 24622
rect 7858 24558 7870 24610
rect 7922 24558 7934 24610
rect 10994 24558 11006 24610
rect 11058 24558 11070 24610
rect 14354 24558 14366 24610
rect 14418 24558 14430 24610
rect 16594 24558 16606 24610
rect 16658 24558 16670 24610
rect 21186 24558 21198 24610
rect 21250 24558 21262 24610
rect 23314 24558 23326 24610
rect 23378 24558 23390 24610
rect 26002 24558 26014 24610
rect 26066 24558 26078 24610
rect 6638 24546 6690 24558
rect 26910 24546 26962 24558
rect 30158 24610 30210 24622
rect 37326 24610 37378 24622
rect 42814 24610 42866 24622
rect 35970 24558 35982 24610
rect 36034 24558 36046 24610
rect 41682 24558 41694 24610
rect 41746 24558 41758 24610
rect 30158 24546 30210 24558
rect 37326 24546 37378 24558
rect 42814 24546 42866 24558
rect 43374 24610 43426 24622
rect 43374 24546 43426 24558
rect 1710 24498 1762 24510
rect 1710 24434 1762 24446
rect 26462 24498 26514 24510
rect 26462 24434 26514 24446
rect 31390 24498 31442 24510
rect 43486 24498 43538 24510
rect 38434 24446 38446 24498
rect 38498 24446 38510 24498
rect 31390 24434 31442 24446
rect 43486 24434 43538 24446
rect 1344 24330 58576 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 58576 24330
rect 1344 24244 58576 24278
rect 5742 24162 5794 24174
rect 46622 24162 46674 24174
rect 19394 24110 19406 24162
rect 19458 24110 19470 24162
rect 5742 24098 5794 24110
rect 46622 24098 46674 24110
rect 46958 24162 47010 24174
rect 46958 24098 47010 24110
rect 47518 24162 47570 24174
rect 47518 24098 47570 24110
rect 5630 24050 5682 24062
rect 20750 24050 20802 24062
rect 31166 24050 31218 24062
rect 6402 23998 6414 24050
rect 6466 23998 6478 24050
rect 18498 23998 18510 24050
rect 18562 23998 18574 24050
rect 19282 23998 19294 24050
rect 19346 23998 19358 24050
rect 28130 23998 28142 24050
rect 28194 23998 28206 24050
rect 5630 23986 5682 23998
rect 20750 23986 20802 23998
rect 31166 23986 31218 23998
rect 40798 24050 40850 24062
rect 45838 24050 45890 24062
rect 43474 23998 43486 24050
rect 43538 23998 43550 24050
rect 40798 23986 40850 23998
rect 45838 23986 45890 23998
rect 46398 24050 46450 24062
rect 46398 23986 46450 23998
rect 57934 24050 57986 24062
rect 57934 23986 57986 23998
rect 14814 23938 14866 23950
rect 15934 23938 15986 23950
rect 22094 23938 22146 23950
rect 22990 23938 23042 23950
rect 27470 23938 27522 23950
rect 29150 23938 29202 23950
rect 41134 23938 41186 23950
rect 7298 23886 7310 23938
rect 7362 23886 7374 23938
rect 8418 23886 8430 23938
rect 8482 23886 8494 23938
rect 9314 23886 9326 23938
rect 9378 23886 9390 23938
rect 9650 23886 9662 23938
rect 9714 23886 9726 23938
rect 10994 23886 11006 23938
rect 11058 23886 11070 23938
rect 11890 23886 11902 23938
rect 11954 23886 11966 23938
rect 14466 23886 14478 23938
rect 14530 23886 14542 23938
rect 15362 23886 15374 23938
rect 15426 23886 15438 23938
rect 16930 23886 16942 23938
rect 16994 23886 17006 23938
rect 17826 23886 17838 23938
rect 17890 23886 17902 23938
rect 18386 23886 18398 23938
rect 18450 23886 18462 23938
rect 19394 23886 19406 23938
rect 19458 23886 19470 23938
rect 22530 23886 22542 23938
rect 22594 23886 22606 23938
rect 24434 23886 24446 23938
rect 24498 23886 24510 23938
rect 26338 23886 26350 23938
rect 26402 23886 26414 23938
rect 28466 23886 28478 23938
rect 28530 23886 28542 23938
rect 29586 23886 29598 23938
rect 29650 23886 29662 23938
rect 31378 23886 31390 23938
rect 31442 23886 31454 23938
rect 33394 23886 33406 23938
rect 33458 23886 33470 23938
rect 14814 23874 14866 23886
rect 15934 23874 15986 23886
rect 22094 23874 22146 23886
rect 22990 23874 23042 23886
rect 27470 23874 27522 23886
rect 29150 23874 29202 23886
rect 41134 23874 41186 23886
rect 41694 23938 41746 23950
rect 42590 23938 42642 23950
rect 47294 23938 47346 23950
rect 42018 23886 42030 23938
rect 42082 23886 42094 23938
rect 43362 23886 43374 23938
rect 43426 23886 43438 23938
rect 55570 23886 55582 23938
rect 55634 23886 55646 23938
rect 41694 23874 41746 23886
rect 42590 23874 42642 23886
rect 47294 23874 47346 23886
rect 34526 23826 34578 23838
rect 9986 23774 9998 23826
rect 10050 23774 10062 23826
rect 11330 23774 11342 23826
rect 11394 23774 11406 23826
rect 12898 23774 12910 23826
rect 12962 23774 12974 23826
rect 15698 23774 15710 23826
rect 15762 23774 15774 23826
rect 16818 23774 16830 23826
rect 16882 23774 16894 23826
rect 23986 23774 23998 23826
rect 24050 23774 24062 23826
rect 26114 23774 26126 23826
rect 26178 23774 26190 23826
rect 31490 23774 31502 23826
rect 31554 23774 31566 23826
rect 34526 23762 34578 23774
rect 44270 23826 44322 23838
rect 44270 23762 44322 23774
rect 45950 23826 46002 23838
rect 50082 23774 50094 23826
rect 50146 23774 50158 23826
rect 45950 23762 46002 23774
rect 13918 23714 13970 23726
rect 21310 23714 21362 23726
rect 40686 23714 40738 23726
rect 17714 23662 17726 23714
rect 17778 23662 17790 23714
rect 25442 23662 25454 23714
rect 25506 23662 25518 23714
rect 27122 23662 27134 23714
rect 27186 23662 27198 23714
rect 35074 23662 35086 23714
rect 35138 23662 35150 23714
rect 13918 23650 13970 23662
rect 21310 23650 21362 23662
rect 40686 23650 40738 23662
rect 42366 23714 42418 23726
rect 42366 23650 42418 23662
rect 42478 23714 42530 23726
rect 42478 23650 42530 23662
rect 45502 23714 45554 23726
rect 45502 23650 45554 23662
rect 45726 23714 45778 23726
rect 49758 23714 49810 23726
rect 47842 23662 47854 23714
rect 47906 23662 47918 23714
rect 45726 23650 45778 23662
rect 49758 23650 49810 23662
rect 1344 23546 58576 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 58576 23546
rect 1344 23460 58576 23494
rect 17614 23378 17666 23390
rect 40910 23378 40962 23390
rect 21858 23326 21870 23378
rect 21922 23326 21934 23378
rect 17614 23314 17666 23326
rect 40910 23314 40962 23326
rect 42590 23378 42642 23390
rect 42590 23314 42642 23326
rect 43150 23378 43202 23390
rect 43150 23314 43202 23326
rect 22430 23266 22482 23278
rect 7746 23214 7758 23266
rect 7810 23214 7822 23266
rect 11666 23214 11678 23266
rect 11730 23214 11742 23266
rect 18834 23214 18846 23266
rect 18898 23214 18910 23266
rect 22430 23202 22482 23214
rect 22654 23266 22706 23278
rect 26014 23266 26066 23278
rect 33742 23266 33794 23278
rect 44942 23266 44994 23278
rect 24658 23214 24670 23266
rect 24722 23214 24734 23266
rect 26338 23214 26350 23266
rect 26402 23214 26414 23266
rect 29474 23214 29486 23266
rect 29538 23214 29550 23266
rect 31378 23214 31390 23266
rect 31442 23214 31454 23266
rect 41234 23214 41246 23266
rect 41298 23214 41310 23266
rect 42802 23214 42814 23266
rect 42866 23214 42878 23266
rect 22654 23202 22706 23214
rect 26014 23202 26066 23214
rect 33742 23202 33794 23214
rect 44942 23202 44994 23214
rect 49758 23266 49810 23278
rect 49758 23202 49810 23214
rect 20638 23154 20690 23166
rect 23102 23154 23154 23166
rect 25678 23154 25730 23166
rect 31950 23154 32002 23166
rect 5058 23102 5070 23154
rect 5122 23102 5134 23154
rect 5618 23102 5630 23154
rect 5682 23102 5694 23154
rect 8418 23102 8430 23154
rect 8482 23102 8494 23154
rect 10210 23102 10222 23154
rect 10274 23102 10286 23154
rect 10994 23102 11006 23154
rect 11058 23102 11070 23154
rect 12786 23102 12798 23154
rect 12850 23102 12862 23154
rect 14130 23102 14142 23154
rect 14194 23102 14206 23154
rect 14914 23102 14926 23154
rect 14978 23102 14990 23154
rect 18050 23102 18062 23154
rect 18114 23102 18126 23154
rect 19618 23102 19630 23154
rect 19682 23102 19694 23154
rect 21410 23102 21422 23154
rect 21474 23102 21486 23154
rect 24322 23102 24334 23154
rect 24386 23102 24398 23154
rect 26674 23102 26686 23154
rect 26738 23102 26750 23154
rect 27458 23102 27470 23154
rect 27522 23102 27534 23154
rect 28242 23102 28254 23154
rect 28306 23102 28318 23154
rect 29922 23102 29934 23154
rect 29986 23102 29998 23154
rect 30930 23102 30942 23154
rect 30994 23102 31006 23154
rect 31266 23102 31278 23154
rect 31330 23102 31342 23154
rect 20638 23090 20690 23102
rect 23102 23090 23154 23102
rect 25678 23090 25730 23102
rect 31950 23090 32002 23102
rect 32510 23154 32562 23166
rect 32510 23090 32562 23102
rect 33518 23154 33570 23166
rect 33518 23090 33570 23102
rect 33630 23154 33682 23166
rect 35758 23154 35810 23166
rect 41918 23154 41970 23166
rect 35074 23102 35086 23154
rect 35138 23102 35150 23154
rect 38882 23102 38894 23154
rect 38946 23102 38958 23154
rect 33630 23090 33682 23102
rect 35758 23090 35810 23102
rect 41918 23090 41970 23102
rect 42142 23154 42194 23166
rect 42142 23090 42194 23102
rect 45390 23154 45442 23166
rect 46162 23102 46174 23154
rect 46226 23102 46238 23154
rect 49074 23102 49086 23154
rect 49138 23102 49150 23154
rect 45390 23090 45442 23102
rect 7198 23042 7250 23054
rect 9998 23042 10050 23054
rect 12238 23042 12290 23054
rect 6514 22990 6526 23042
rect 6578 22990 6590 23042
rect 7746 22990 7758 23042
rect 7810 22990 7822 23042
rect 10882 22990 10894 23042
rect 10946 22990 10958 23042
rect 7198 22978 7250 22990
rect 9998 22978 10050 22990
rect 12238 22978 12290 22990
rect 15710 23042 15762 23054
rect 15710 22978 15762 22990
rect 16158 23042 16210 23054
rect 16158 22978 16210 22990
rect 16606 23042 16658 23054
rect 34302 23042 34354 23054
rect 38334 23042 38386 23054
rect 41694 23042 41746 23054
rect 22754 22990 22766 23042
rect 22818 22990 22830 23042
rect 24434 22990 24446 23042
rect 24498 22990 24510 23042
rect 25330 22990 25342 23042
rect 25394 22990 25406 23042
rect 26898 22990 26910 23042
rect 26962 22990 26974 23042
rect 29026 22990 29038 23042
rect 29090 22990 29102 23042
rect 34850 22990 34862 23042
rect 34914 22990 34926 23042
rect 39106 22990 39118 23042
rect 39170 22990 39182 23042
rect 16606 22978 16658 22990
rect 34302 22978 34354 22990
rect 38334 22978 38386 22990
rect 41694 22978 41746 22990
rect 44606 23042 44658 23054
rect 46846 23042 46898 23054
rect 46386 22990 46398 23042
rect 46450 22990 46462 23042
rect 48850 22990 48862 23042
rect 48914 22990 48926 23042
rect 44606 22978 44658 22990
rect 46846 22978 46898 22990
rect 23326 22930 23378 22942
rect 45054 22930 45106 22942
rect 13906 22878 13918 22930
rect 13970 22878 13982 22930
rect 15474 22878 15486 22930
rect 15538 22927 15550 22930
rect 16370 22927 16382 22930
rect 15538 22881 16382 22927
rect 15538 22878 15550 22881
rect 16370 22878 16382 22881
rect 16434 22878 16446 22930
rect 23650 22878 23662 22930
rect 23714 22878 23726 22930
rect 33058 22878 33070 22930
rect 33122 22878 33134 22930
rect 39330 22878 39342 22930
rect 39394 22878 39406 22930
rect 23326 22866 23378 22878
rect 45054 22866 45106 22878
rect 45502 22930 45554 22942
rect 45502 22866 45554 22878
rect 1344 22762 58576 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 58576 22762
rect 1344 22676 58576 22710
rect 26574 22594 26626 22606
rect 45614 22594 45666 22606
rect 29138 22542 29150 22594
rect 29202 22591 29214 22594
rect 29202 22545 29423 22591
rect 29202 22542 29214 22545
rect 26574 22530 26626 22542
rect 10110 22482 10162 22494
rect 10110 22418 10162 22430
rect 16718 22482 16770 22494
rect 20302 22482 20354 22494
rect 17602 22430 17614 22482
rect 17666 22430 17678 22482
rect 16718 22418 16770 22430
rect 20302 22418 20354 22430
rect 20750 22482 20802 22494
rect 20750 22418 20802 22430
rect 25454 22482 25506 22494
rect 29377 22479 29423 22545
rect 45614 22530 45666 22542
rect 49198 22594 49250 22606
rect 49198 22530 49250 22542
rect 31502 22482 31554 22494
rect 38334 22482 38386 22494
rect 48974 22482 49026 22494
rect 29810 22479 29822 22482
rect 29377 22433 29822 22479
rect 29810 22430 29822 22433
rect 29874 22430 29886 22482
rect 33394 22430 33406 22482
rect 33458 22430 33470 22482
rect 35186 22430 35198 22482
rect 35250 22430 35262 22482
rect 36194 22430 36206 22482
rect 36258 22430 36270 22482
rect 37762 22430 37774 22482
rect 37826 22430 37838 22482
rect 39218 22430 39230 22482
rect 39282 22430 39294 22482
rect 40450 22430 40462 22482
rect 40514 22430 40526 22482
rect 25454 22418 25506 22430
rect 31502 22418 31554 22430
rect 38334 22418 38386 22430
rect 48974 22418 49026 22430
rect 57934 22482 57986 22494
rect 57934 22418 57986 22430
rect 6078 22370 6130 22382
rect 6078 22306 6130 22318
rect 6638 22370 6690 22382
rect 6638 22306 6690 22318
rect 6974 22370 7026 22382
rect 8990 22370 9042 22382
rect 25902 22370 25954 22382
rect 8530 22318 8542 22370
rect 8594 22318 8606 22370
rect 10546 22318 10558 22370
rect 10610 22318 10622 22370
rect 12450 22318 12462 22370
rect 12514 22318 12526 22370
rect 14130 22318 14142 22370
rect 14194 22318 14206 22370
rect 15810 22318 15822 22370
rect 15874 22318 15886 22370
rect 16258 22318 16270 22370
rect 16322 22318 16334 22370
rect 17266 22318 17278 22370
rect 17330 22318 17342 22370
rect 18050 22318 18062 22370
rect 18114 22318 18126 22370
rect 19170 22318 19182 22370
rect 19234 22318 19246 22370
rect 19730 22318 19742 22370
rect 19794 22318 19806 22370
rect 20178 22318 20190 22370
rect 20242 22318 20254 22370
rect 21410 22318 21422 22370
rect 21474 22318 21486 22370
rect 21634 22318 21646 22370
rect 21698 22318 21710 22370
rect 23538 22318 23550 22370
rect 23602 22318 23614 22370
rect 6974 22306 7026 22318
rect 8990 22306 9042 22318
rect 25902 22306 25954 22318
rect 26126 22370 26178 22382
rect 26126 22306 26178 22318
rect 26462 22370 26514 22382
rect 26462 22306 26514 22318
rect 26686 22370 26738 22382
rect 26686 22306 26738 22318
rect 27022 22370 27074 22382
rect 27022 22306 27074 22318
rect 27582 22370 27634 22382
rect 35758 22370 35810 22382
rect 40014 22370 40066 22382
rect 28466 22318 28478 22370
rect 28530 22318 28542 22370
rect 29810 22318 29822 22370
rect 29874 22318 29886 22370
rect 31938 22318 31950 22370
rect 32002 22318 32014 22370
rect 33842 22318 33854 22370
rect 33906 22318 33918 22370
rect 34962 22318 34974 22370
rect 35026 22318 35038 22370
rect 35970 22318 35982 22370
rect 36034 22318 36046 22370
rect 38994 22318 39006 22370
rect 39058 22318 39070 22370
rect 27582 22306 27634 22318
rect 35758 22306 35810 22318
rect 40014 22306 40066 22318
rect 44942 22370 44994 22382
rect 45726 22370 45778 22382
rect 45266 22318 45278 22370
rect 45330 22318 45342 22370
rect 44942 22306 44994 22318
rect 45726 22306 45778 22318
rect 46398 22370 46450 22382
rect 55570 22318 55582 22370
rect 55634 22318 55646 22370
rect 46398 22306 46450 22318
rect 7534 22258 7586 22270
rect 12014 22258 12066 22270
rect 28030 22258 28082 22270
rect 11554 22206 11566 22258
rect 11618 22206 11630 22258
rect 13458 22206 13470 22258
rect 13522 22206 13534 22258
rect 18162 22206 18174 22258
rect 18226 22206 18238 22258
rect 24658 22206 24670 22258
rect 24722 22206 24734 22258
rect 7534 22194 7586 22206
rect 12014 22194 12066 22206
rect 28030 22194 28082 22206
rect 29262 22258 29314 22270
rect 37214 22258 37266 22270
rect 30930 22206 30942 22258
rect 30994 22206 31006 22258
rect 32386 22206 32398 22258
rect 32450 22206 32462 22258
rect 29262 22194 29314 22206
rect 37214 22194 37266 22206
rect 37326 22258 37378 22270
rect 39678 22258 39730 22270
rect 37426 22206 37438 22258
rect 37490 22206 37502 22258
rect 37326 22194 37378 22206
rect 39678 22194 39730 22206
rect 46174 22258 46226 22270
rect 46174 22194 46226 22206
rect 8094 22146 8146 22158
rect 15710 22146 15762 22158
rect 24894 22146 24946 22158
rect 8306 22094 8318 22146
rect 8370 22094 8382 22146
rect 9314 22094 9326 22146
rect 9378 22094 9390 22146
rect 18946 22094 18958 22146
rect 19010 22094 19022 22146
rect 8094 22082 8146 22094
rect 15710 22082 15762 22094
rect 24894 22082 24946 22094
rect 36990 22146 37042 22158
rect 36990 22082 37042 22094
rect 45502 22146 45554 22158
rect 45502 22082 45554 22094
rect 46286 22146 46338 22158
rect 49522 22094 49534 22146
rect 49586 22094 49598 22146
rect 46286 22082 46338 22094
rect 1344 21978 58576 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 58576 21978
rect 1344 21892 58576 21926
rect 5630 21810 5682 21822
rect 5630 21746 5682 21758
rect 5854 21810 5906 21822
rect 5854 21746 5906 21758
rect 10334 21810 10386 21822
rect 10334 21746 10386 21758
rect 17726 21810 17778 21822
rect 17726 21746 17778 21758
rect 22430 21810 22482 21822
rect 22430 21746 22482 21758
rect 26014 21810 26066 21822
rect 26014 21746 26066 21758
rect 26798 21810 26850 21822
rect 26798 21746 26850 21758
rect 27806 21810 27858 21822
rect 27806 21746 27858 21758
rect 28366 21810 28418 21822
rect 32062 21810 32114 21822
rect 29586 21758 29598 21810
rect 29650 21758 29662 21810
rect 28366 21746 28418 21758
rect 32062 21746 32114 21758
rect 33854 21810 33906 21822
rect 41694 21810 41746 21822
rect 35186 21758 35198 21810
rect 35250 21758 35262 21810
rect 33854 21746 33906 21758
rect 41694 21746 41746 21758
rect 42142 21810 42194 21822
rect 58158 21810 58210 21822
rect 42466 21758 42478 21810
rect 42530 21758 42542 21810
rect 51090 21758 51102 21810
rect 51154 21758 51166 21810
rect 42142 21746 42194 21758
rect 58158 21746 58210 21758
rect 1710 21698 1762 21710
rect 14254 21698 14306 21710
rect 26238 21698 26290 21710
rect 31054 21698 31106 21710
rect 11554 21646 11566 21698
rect 11618 21646 11630 21698
rect 20178 21646 20190 21698
rect 20242 21646 20254 21698
rect 21186 21646 21198 21698
rect 21250 21646 21262 21698
rect 28914 21646 28926 21698
rect 28978 21646 28990 21698
rect 29138 21646 29150 21698
rect 29202 21646 29214 21698
rect 1710 21634 1762 21646
rect 14254 21634 14306 21646
rect 26238 21634 26290 21646
rect 31054 21634 31106 21646
rect 31166 21698 31218 21710
rect 31166 21634 31218 21646
rect 32398 21698 32450 21710
rect 37550 21698 37602 21710
rect 35074 21646 35086 21698
rect 35138 21646 35150 21698
rect 32398 21634 32450 21646
rect 37550 21634 37602 21646
rect 42814 21698 42866 21710
rect 42814 21634 42866 21646
rect 43038 21698 43090 21710
rect 43038 21634 43090 21646
rect 43374 21698 43426 21710
rect 43374 21634 43426 21646
rect 6414 21586 6466 21598
rect 16158 21586 16210 21598
rect 7298 21534 7310 21586
rect 7362 21534 7374 21586
rect 11218 21534 11230 21586
rect 11282 21534 11294 21586
rect 14802 21534 14814 21586
rect 14866 21534 14878 21586
rect 6414 21522 6466 21534
rect 16158 21522 16210 21534
rect 18622 21586 18674 21598
rect 23438 21586 23490 21598
rect 25230 21586 25282 21598
rect 19058 21534 19070 21586
rect 19122 21534 19134 21586
rect 20290 21534 20302 21586
rect 20354 21534 20366 21586
rect 21074 21534 21086 21586
rect 21138 21534 21150 21586
rect 21858 21534 21870 21586
rect 21922 21534 21934 21586
rect 23090 21534 23102 21586
rect 23154 21534 23166 21586
rect 24322 21534 24334 21586
rect 24386 21534 24398 21586
rect 18622 21522 18674 21534
rect 23438 21522 23490 21534
rect 25230 21522 25282 21534
rect 25342 21586 25394 21598
rect 25342 21522 25394 21534
rect 25454 21586 25506 21598
rect 26350 21586 26402 21598
rect 30046 21586 30098 21598
rect 25778 21534 25790 21586
rect 25842 21534 25854 21586
rect 28578 21534 28590 21586
rect 28642 21534 28654 21586
rect 25454 21522 25506 21534
rect 26350 21522 26402 21534
rect 30046 21522 30098 21534
rect 30830 21586 30882 21598
rect 30830 21522 30882 21534
rect 33070 21586 33122 21598
rect 33070 21522 33122 21534
rect 33294 21586 33346 21598
rect 33294 21522 33346 21534
rect 33518 21586 33570 21598
rect 33518 21522 33570 21534
rect 33742 21586 33794 21598
rect 33742 21522 33794 21534
rect 34078 21586 34130 21598
rect 38670 21586 38722 21598
rect 41582 21586 41634 21598
rect 50430 21586 50482 21598
rect 34962 21534 34974 21586
rect 35026 21534 35038 21586
rect 39554 21534 39566 21586
rect 39618 21534 39630 21586
rect 49746 21534 49758 21586
rect 49810 21534 49822 21586
rect 34078 21522 34130 21534
rect 38670 21522 38722 21534
rect 41582 21522 41634 21534
rect 50430 21522 50482 21534
rect 50766 21586 50818 21598
rect 50766 21522 50818 21534
rect 6974 21474 7026 21486
rect 8990 21474 9042 21486
rect 7970 21422 7982 21474
rect 8034 21422 8046 21474
rect 6974 21410 7026 21422
rect 8990 21410 9042 21422
rect 10110 21474 10162 21486
rect 10110 21410 10162 21422
rect 10894 21474 10946 21486
rect 12462 21474 12514 21486
rect 11890 21422 11902 21474
rect 11954 21422 11966 21474
rect 10894 21410 10946 21422
rect 12462 21410 12514 21422
rect 12910 21474 12962 21486
rect 12910 21410 12962 21422
rect 15038 21474 15090 21486
rect 15038 21410 15090 21422
rect 15598 21474 15650 21486
rect 18286 21474 18338 21486
rect 16594 21422 16606 21474
rect 16658 21422 16670 21474
rect 15598 21410 15650 21422
rect 18286 21410 18338 21422
rect 19854 21474 19906 21486
rect 27246 21474 27298 21486
rect 23874 21422 23886 21474
rect 23938 21422 23950 21474
rect 19854 21410 19906 21422
rect 27246 21410 27298 21422
rect 30606 21474 30658 21486
rect 30606 21410 30658 21422
rect 31726 21474 31778 21486
rect 31726 21410 31778 21422
rect 34638 21474 34690 21486
rect 43262 21474 43314 21486
rect 39218 21422 39230 21474
rect 39282 21422 39294 21474
rect 49522 21422 49534 21474
rect 49586 21422 49598 21474
rect 34638 21410 34690 21422
rect 43262 21410 43314 21422
rect 32510 21362 32562 21374
rect 24210 21310 24222 21362
rect 24274 21310 24286 21362
rect 32510 21298 32562 21310
rect 41694 21362 41746 21374
rect 41694 21298 41746 21310
rect 1344 21194 58576 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 58576 21194
rect 1344 21108 58576 21142
rect 17054 21026 17106 21038
rect 35646 21026 35698 21038
rect 31826 20974 31838 21026
rect 31890 20974 31902 21026
rect 33842 20974 33854 21026
rect 33906 20974 33918 21026
rect 17054 20962 17106 20974
rect 35646 20962 35698 20974
rect 8990 20914 9042 20926
rect 18174 20914 18226 20926
rect 6962 20862 6974 20914
rect 7026 20862 7038 20914
rect 11330 20862 11342 20914
rect 11394 20862 11406 20914
rect 12226 20862 12238 20914
rect 12290 20862 12302 20914
rect 13906 20862 13918 20914
rect 13970 20862 13982 20914
rect 16706 20862 16718 20914
rect 16770 20862 16782 20914
rect 8990 20850 9042 20862
rect 18174 20850 18226 20862
rect 35870 20914 35922 20926
rect 35870 20850 35922 20862
rect 36206 20914 36258 20926
rect 36206 20850 36258 20862
rect 37662 20914 37714 20926
rect 37662 20850 37714 20862
rect 38670 20914 38722 20926
rect 38670 20850 38722 20862
rect 42366 20914 42418 20926
rect 42366 20850 42418 20862
rect 43710 20914 43762 20926
rect 43710 20850 43762 20862
rect 44046 20914 44098 20926
rect 44046 20850 44098 20862
rect 48638 20914 48690 20926
rect 49522 20862 49534 20914
rect 49586 20862 49598 20914
rect 48638 20850 48690 20862
rect 8094 20802 8146 20814
rect 11790 20802 11842 20814
rect 16270 20802 16322 20814
rect 7522 20750 7534 20802
rect 7586 20750 7598 20802
rect 10210 20750 10222 20802
rect 10274 20750 10286 20802
rect 13682 20750 13694 20802
rect 13746 20750 13758 20802
rect 15810 20750 15822 20802
rect 15874 20750 15886 20802
rect 8094 20738 8146 20750
rect 11790 20738 11842 20750
rect 16270 20738 16322 20750
rect 16494 20802 16546 20814
rect 16494 20738 16546 20750
rect 17390 20802 17442 20814
rect 28030 20802 28082 20814
rect 33518 20802 33570 20814
rect 17602 20750 17614 20802
rect 17666 20750 17678 20802
rect 19394 20750 19406 20802
rect 19458 20750 19470 20802
rect 22194 20750 22206 20802
rect 22258 20750 22270 20802
rect 23762 20750 23774 20802
rect 23826 20750 23838 20802
rect 25330 20750 25342 20802
rect 25394 20750 25406 20802
rect 26226 20750 26238 20802
rect 26290 20750 26302 20802
rect 27234 20750 27246 20802
rect 27298 20750 27310 20802
rect 28466 20750 28478 20802
rect 28530 20750 28542 20802
rect 29586 20750 29598 20802
rect 29650 20750 29662 20802
rect 30706 20750 30718 20802
rect 30770 20750 30782 20802
rect 31602 20750 31614 20802
rect 31666 20750 31678 20802
rect 17390 20738 17442 20750
rect 28030 20738 28082 20750
rect 33518 20738 33570 20750
rect 34638 20802 34690 20814
rect 34638 20738 34690 20750
rect 35086 20802 35138 20814
rect 35086 20738 35138 20750
rect 36318 20802 36370 20814
rect 41134 20802 41186 20814
rect 41582 20802 41634 20814
rect 42814 20802 42866 20814
rect 38098 20750 38110 20802
rect 38162 20750 38174 20802
rect 39666 20750 39678 20802
rect 39730 20750 39742 20802
rect 41346 20750 41358 20802
rect 41410 20750 41422 20802
rect 41682 20750 41694 20802
rect 41746 20750 41758 20802
rect 43250 20750 43262 20802
rect 43314 20750 43326 20802
rect 47282 20750 47294 20802
rect 47346 20750 47358 20802
rect 47954 20750 47966 20802
rect 48018 20750 48030 20802
rect 48850 20750 48862 20802
rect 48914 20750 48926 20802
rect 49746 20750 49758 20802
rect 49810 20750 49822 20802
rect 36318 20738 36370 20750
rect 41134 20738 41186 20750
rect 41582 20738 41634 20750
rect 42814 20738 42866 20750
rect 6302 20690 6354 20702
rect 6302 20626 6354 20638
rect 8654 20690 8706 20702
rect 8654 20626 8706 20638
rect 12686 20690 12738 20702
rect 16830 20690 16882 20702
rect 26014 20690 26066 20702
rect 27022 20690 27074 20702
rect 34974 20690 35026 20702
rect 40910 20690 40962 20702
rect 13458 20638 13470 20690
rect 13522 20638 13534 20690
rect 19282 20638 19294 20690
rect 19346 20638 19358 20690
rect 22306 20638 22318 20690
rect 22370 20638 22382 20690
rect 26786 20638 26798 20690
rect 26850 20638 26862 20690
rect 31938 20638 31950 20690
rect 32002 20638 32014 20690
rect 39890 20638 39902 20690
rect 39954 20638 39966 20690
rect 40338 20638 40350 20690
rect 40402 20638 40414 20690
rect 12686 20626 12738 20638
rect 16830 20626 16882 20638
rect 26014 20626 26066 20638
rect 27022 20626 27074 20638
rect 34974 20626 35026 20638
rect 40910 20626 40962 20638
rect 45614 20690 45666 20702
rect 45614 20626 45666 20638
rect 46062 20690 46114 20702
rect 46062 20626 46114 20638
rect 46174 20690 46226 20702
rect 46722 20638 46734 20690
rect 46786 20638 46798 20690
rect 50306 20638 50318 20690
rect 50370 20638 50382 20690
rect 46174 20626 46226 20638
rect 9550 20578 9602 20590
rect 9550 20514 9602 20526
rect 12798 20578 12850 20590
rect 12798 20514 12850 20526
rect 13022 20578 13074 20590
rect 13022 20514 13074 20526
rect 18622 20578 18674 20590
rect 21646 20578 21698 20590
rect 36094 20578 36146 20590
rect 20626 20526 20638 20578
rect 20690 20526 20702 20578
rect 22418 20526 22430 20578
rect 22482 20526 22494 20578
rect 18622 20514 18674 20526
rect 21646 20514 21698 20526
rect 36094 20514 36146 20526
rect 41918 20578 41970 20590
rect 41918 20514 41970 20526
rect 44158 20578 44210 20590
rect 44158 20514 44210 20526
rect 45838 20578 45890 20590
rect 45838 20514 45890 20526
rect 1344 20410 58576 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 58576 20410
rect 1344 20324 58576 20358
rect 22094 20242 22146 20254
rect 30718 20242 30770 20254
rect 16594 20190 16606 20242
rect 16658 20190 16670 20242
rect 18946 20190 18958 20242
rect 19010 20190 19022 20242
rect 23314 20190 23326 20242
rect 23378 20190 23390 20242
rect 22094 20178 22146 20190
rect 30718 20178 30770 20190
rect 31726 20242 31778 20254
rect 31726 20178 31778 20190
rect 31838 20242 31890 20254
rect 31838 20178 31890 20190
rect 34862 20242 34914 20254
rect 58158 20242 58210 20254
rect 40226 20190 40238 20242
rect 40290 20190 40302 20242
rect 34862 20178 34914 20190
rect 58158 20178 58210 20190
rect 5294 20130 5346 20142
rect 18062 20130 18114 20142
rect 24222 20130 24274 20142
rect 26574 20130 26626 20142
rect 9762 20078 9774 20130
rect 9826 20078 9838 20130
rect 15138 20078 15150 20130
rect 15202 20078 15214 20130
rect 19170 20078 19182 20130
rect 19234 20078 19246 20130
rect 19730 20078 19742 20130
rect 19794 20078 19806 20130
rect 22418 20078 22430 20130
rect 22482 20078 22494 20130
rect 25554 20078 25566 20130
rect 25618 20078 25630 20130
rect 5294 20066 5346 20078
rect 18062 20066 18114 20078
rect 24222 20066 24274 20078
rect 26574 20066 26626 20078
rect 27470 20130 27522 20142
rect 49198 20130 49250 20142
rect 28130 20078 28142 20130
rect 28194 20078 28206 20130
rect 28578 20078 28590 20130
rect 28642 20078 28654 20130
rect 33282 20078 33294 20130
rect 33346 20078 33358 20130
rect 33618 20078 33630 20130
rect 33682 20078 33694 20130
rect 34514 20078 34526 20130
rect 34578 20078 34590 20130
rect 36194 20078 36206 20130
rect 36258 20078 36270 20130
rect 39442 20078 39454 20130
rect 39506 20078 39518 20130
rect 41570 20078 41582 20130
rect 41634 20078 41646 20130
rect 46162 20078 46174 20130
rect 46226 20078 46238 20130
rect 46722 20078 46734 20130
rect 46786 20078 46798 20130
rect 27470 20066 27522 20078
rect 49198 20066 49250 20078
rect 49310 20130 49362 20142
rect 49310 20066 49362 20078
rect 5854 20018 5906 20030
rect 19406 20018 19458 20030
rect 23998 20018 24050 20030
rect 7074 19966 7086 20018
rect 7138 19966 7150 20018
rect 8530 19966 8542 20018
rect 8594 19966 8606 20018
rect 9538 19966 9550 20018
rect 9602 19966 9614 20018
rect 10882 19966 10894 20018
rect 10946 19966 10958 20018
rect 12450 19966 12462 20018
rect 12514 19966 12526 20018
rect 13010 19966 13022 20018
rect 13074 19966 13086 20018
rect 13458 19966 13470 20018
rect 13522 19966 13534 20018
rect 13682 19966 13694 20018
rect 13746 19966 13758 20018
rect 16594 19966 16606 20018
rect 16658 19966 16670 20018
rect 18610 19966 18622 20018
rect 18674 19966 18686 20018
rect 20066 19966 20078 20018
rect 20130 19966 20142 20018
rect 21074 19966 21086 20018
rect 21138 19966 21150 20018
rect 21298 19966 21310 20018
rect 21362 19966 21374 20018
rect 22306 19966 22318 20018
rect 22370 19966 22382 20018
rect 23426 19966 23438 20018
rect 23490 19966 23502 20018
rect 5854 19954 5906 19966
rect 19406 19954 19458 19966
rect 23998 19954 24050 19966
rect 24446 20018 24498 20030
rect 24446 19954 24498 19966
rect 24558 20018 24610 20030
rect 27582 20018 27634 20030
rect 25330 19966 25342 20018
rect 25394 19966 25406 20018
rect 26226 19966 26238 20018
rect 26290 19966 26302 20018
rect 24558 19954 24610 19966
rect 27582 19954 27634 19966
rect 27694 20018 27746 20030
rect 31614 20018 31666 20030
rect 28802 19966 28814 20018
rect 28866 19966 28878 20018
rect 30818 19966 30830 20018
rect 30882 19966 30894 20018
rect 27694 19954 27746 19966
rect 31614 19954 31666 19966
rect 31950 20018 32002 20030
rect 36542 20018 36594 20030
rect 32162 19966 32174 20018
rect 32226 19966 32238 20018
rect 33058 19966 33070 20018
rect 33122 19966 33134 20018
rect 35970 19966 35982 20018
rect 36034 19966 36046 20018
rect 31950 19954 32002 19966
rect 36542 19954 36594 19966
rect 37886 20018 37938 20030
rect 37886 19954 37938 19966
rect 38334 20018 38386 20030
rect 38334 19954 38386 19966
rect 38558 20018 38610 20030
rect 42702 20018 42754 20030
rect 44718 20018 44770 20030
rect 49534 20018 49586 20030
rect 39330 19966 39342 20018
rect 39394 19966 39406 20018
rect 40114 19966 40126 20018
rect 40178 19966 40190 20018
rect 41906 19966 41918 20018
rect 41970 19966 41982 20018
rect 42914 19966 42926 20018
rect 42978 19966 42990 20018
rect 44930 19966 44942 20018
rect 44994 19966 45006 20018
rect 46050 19966 46062 20018
rect 46114 19966 46126 20018
rect 46834 19966 46846 20018
rect 46898 19966 46910 20018
rect 47506 19966 47518 20018
rect 47570 19966 47582 20018
rect 47954 19966 47966 20018
rect 48018 19966 48030 20018
rect 38558 19954 38610 19966
rect 42702 19954 42754 19966
rect 44718 19954 44770 19966
rect 49534 19954 49586 19966
rect 4958 19906 5010 19918
rect 11342 19906 11394 19918
rect 34302 19906 34354 19918
rect 7410 19854 7422 19906
rect 7474 19903 7486 19906
rect 7634 19903 7646 19906
rect 7474 19857 7646 19903
rect 7474 19854 7486 19857
rect 7634 19854 7646 19857
rect 7698 19854 7710 19906
rect 8418 19854 8430 19906
rect 8482 19854 8494 19906
rect 10210 19854 10222 19906
rect 10274 19854 10286 19906
rect 17602 19854 17614 19906
rect 17666 19854 17678 19906
rect 20402 19854 20414 19906
rect 20466 19854 20478 19906
rect 20850 19854 20862 19906
rect 20914 19854 20926 19906
rect 26002 19854 26014 19906
rect 26066 19854 26078 19906
rect 4958 19842 5010 19854
rect 11342 19842 11394 19854
rect 34302 19842 34354 19854
rect 37102 19906 37154 19918
rect 37102 19842 37154 19854
rect 38446 19906 38498 19918
rect 45938 19854 45950 19906
rect 46002 19854 46014 19906
rect 38446 19842 38498 19854
rect 18958 19794 19010 19806
rect 8754 19742 8766 19794
rect 8818 19742 8830 19794
rect 43698 19742 43710 19794
rect 43762 19742 43774 19794
rect 47058 19742 47070 19794
rect 47122 19742 47134 19794
rect 18958 19730 19010 19742
rect 1344 19626 58576 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 58576 19626
rect 1344 19540 58576 19574
rect 6750 19458 6802 19470
rect 6750 19394 6802 19406
rect 17502 19458 17554 19470
rect 17502 19394 17554 19406
rect 17838 19458 17890 19470
rect 17838 19394 17890 19406
rect 23886 19458 23938 19470
rect 23886 19394 23938 19406
rect 23998 19458 24050 19470
rect 23998 19394 24050 19406
rect 24222 19458 24274 19470
rect 43710 19458 43762 19470
rect 40674 19406 40686 19458
rect 40738 19406 40750 19458
rect 24222 19394 24274 19406
rect 43710 19394 43762 19406
rect 44270 19458 44322 19470
rect 44270 19394 44322 19406
rect 46958 19458 47010 19470
rect 46958 19394 47010 19406
rect 49198 19458 49250 19470
rect 49198 19394 49250 19406
rect 13582 19346 13634 19358
rect 11554 19294 11566 19346
rect 11618 19294 11630 19346
rect 13582 19282 13634 19294
rect 14142 19346 14194 19358
rect 18398 19346 18450 19358
rect 25118 19346 25170 19358
rect 15026 19294 15038 19346
rect 15090 19294 15102 19346
rect 21410 19294 21422 19346
rect 21474 19294 21486 19346
rect 14142 19282 14194 19294
rect 18398 19282 18450 19294
rect 25118 19282 25170 19294
rect 27582 19346 27634 19358
rect 27582 19282 27634 19294
rect 28142 19346 28194 19358
rect 28142 19282 28194 19294
rect 32734 19346 32786 19358
rect 48974 19346 49026 19358
rect 38210 19294 38222 19346
rect 38274 19294 38286 19346
rect 44034 19294 44046 19346
rect 44098 19294 44110 19346
rect 32734 19282 32786 19294
rect 48974 19282 49026 19294
rect 50094 19346 50146 19358
rect 50094 19282 50146 19294
rect 5630 19234 5682 19246
rect 5630 19170 5682 19182
rect 6526 19234 6578 19246
rect 6526 19170 6578 19182
rect 7646 19234 7698 19246
rect 7646 19170 7698 19182
rect 7870 19234 7922 19246
rect 7870 19170 7922 19182
rect 8318 19234 8370 19246
rect 8318 19170 8370 19182
rect 9102 19234 9154 19246
rect 9102 19170 9154 19182
rect 9662 19234 9714 19246
rect 18734 19234 18786 19246
rect 11442 19182 11454 19234
rect 11506 19182 11518 19234
rect 12002 19182 12014 19234
rect 12066 19182 12078 19234
rect 14242 19182 14254 19234
rect 14306 19182 14318 19234
rect 15250 19182 15262 19234
rect 15314 19182 15326 19234
rect 15922 19182 15934 19234
rect 15986 19182 15998 19234
rect 9662 19170 9714 19182
rect 18734 19170 18786 19182
rect 19182 19234 19234 19246
rect 22766 19234 22818 19246
rect 20290 19182 20302 19234
rect 20354 19182 20366 19234
rect 21858 19182 21870 19234
rect 21922 19182 21934 19234
rect 19182 19170 19234 19182
rect 22766 19170 22818 19182
rect 22990 19234 23042 19246
rect 22990 19170 23042 19182
rect 25678 19234 25730 19246
rect 26238 19234 26290 19246
rect 26002 19182 26014 19234
rect 26066 19182 26078 19234
rect 25678 19170 25730 19182
rect 26238 19170 26290 19182
rect 29262 19234 29314 19246
rect 29262 19170 29314 19182
rect 29598 19234 29650 19246
rect 29598 19170 29650 19182
rect 29934 19234 29986 19246
rect 29934 19170 29986 19182
rect 36430 19234 36482 19246
rect 40014 19234 40066 19246
rect 37426 19182 37438 19234
rect 37490 19182 37502 19234
rect 38322 19182 38334 19234
rect 38386 19182 38398 19234
rect 36430 19170 36482 19182
rect 40014 19170 40066 19182
rect 43486 19234 43538 19246
rect 43486 19170 43538 19182
rect 46286 19234 46338 19246
rect 46610 19182 46622 19234
rect 46674 19182 46686 19234
rect 51426 19182 51438 19234
rect 51490 19182 51502 19234
rect 46286 19170 46338 19182
rect 7086 19122 7138 19134
rect 22318 19122 22370 19134
rect 10882 19070 10894 19122
rect 10946 19070 10958 19122
rect 15698 19070 15710 19122
rect 15762 19070 15774 19122
rect 16258 19070 16270 19122
rect 16322 19070 16334 19122
rect 16930 19070 16942 19122
rect 16994 19070 17006 19122
rect 17266 19070 17278 19122
rect 17330 19070 17342 19122
rect 19954 19070 19966 19122
rect 20018 19070 20030 19122
rect 7086 19058 7138 19070
rect 22318 19058 22370 19070
rect 22878 19122 22930 19134
rect 22878 19058 22930 19070
rect 25902 19122 25954 19134
rect 25902 19058 25954 19070
rect 37214 19122 37266 19134
rect 40126 19122 40178 19134
rect 38546 19070 38558 19122
rect 38610 19070 38622 19122
rect 37214 19058 37266 19070
rect 40126 19058 40178 19070
rect 40238 19122 40290 19134
rect 40238 19058 40290 19070
rect 44046 19122 44098 19134
rect 52110 19122 52162 19134
rect 49522 19070 49534 19122
rect 49586 19070 49598 19122
rect 50194 19070 50206 19122
rect 50258 19070 50270 19122
rect 44046 19058 44098 19070
rect 52110 19058 52162 19070
rect 52670 19122 52722 19134
rect 52670 19058 52722 19070
rect 7758 19010 7810 19022
rect 5954 18958 5966 19010
rect 6018 18958 6030 19010
rect 7758 18946 7810 18958
rect 8990 19010 9042 19022
rect 8990 18946 9042 18958
rect 9550 19010 9602 19022
rect 9550 18946 9602 18958
rect 9774 19010 9826 19022
rect 9774 18946 9826 18958
rect 18846 19010 18898 19022
rect 23886 19010 23938 19022
rect 20402 18958 20414 19010
rect 20466 18958 20478 19010
rect 23426 18958 23438 19010
rect 23490 18958 23502 19010
rect 18846 18946 18898 18958
rect 23886 18946 23938 18958
rect 25006 19010 25058 19022
rect 25006 18946 25058 18958
rect 25230 19010 25282 19022
rect 25230 18946 25282 18958
rect 27134 19010 27186 19022
rect 27134 18946 27186 18958
rect 28590 19010 28642 19022
rect 28590 18946 28642 18958
rect 29598 19010 29650 19022
rect 29598 18946 29650 18958
rect 30382 19010 30434 19022
rect 30382 18946 30434 18958
rect 31166 19010 31218 19022
rect 31166 18946 31218 18958
rect 31614 19010 31666 19022
rect 33966 19010 34018 19022
rect 33618 18958 33630 19010
rect 33682 18958 33694 19010
rect 31614 18946 31666 18958
rect 33966 18946 34018 18958
rect 35870 19010 35922 19022
rect 35870 18946 35922 18958
rect 42366 19010 42418 19022
rect 42366 18946 42418 18958
rect 46846 19010 46898 19022
rect 46846 18946 46898 18958
rect 53006 19010 53058 19022
rect 53006 18946 53058 18958
rect 58158 19010 58210 19022
rect 58158 18946 58210 18958
rect 1344 18842 58576 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 58576 18842
rect 1344 18756 58576 18790
rect 7310 18674 7362 18686
rect 24670 18674 24722 18686
rect 11330 18622 11342 18674
rect 11394 18622 11406 18674
rect 19394 18622 19406 18674
rect 19458 18622 19470 18674
rect 24210 18622 24222 18674
rect 24274 18671 24286 18674
rect 24434 18671 24446 18674
rect 24274 18625 24446 18671
rect 24274 18622 24286 18625
rect 24434 18622 24446 18625
rect 24498 18622 24510 18674
rect 7310 18610 7362 18622
rect 24670 18610 24722 18622
rect 26686 18674 26738 18686
rect 26686 18610 26738 18622
rect 28478 18674 28530 18686
rect 43586 18622 43598 18674
rect 43650 18622 43662 18674
rect 28478 18610 28530 18622
rect 5182 18562 5234 18574
rect 5182 18498 5234 18510
rect 7198 18562 7250 18574
rect 8990 18562 9042 18574
rect 16718 18562 16770 18574
rect 7970 18510 7982 18562
rect 8034 18510 8046 18562
rect 8306 18510 8318 18562
rect 8370 18510 8382 18562
rect 10322 18510 10334 18562
rect 10386 18510 10398 18562
rect 15810 18510 15822 18562
rect 15874 18510 15886 18562
rect 16258 18510 16270 18562
rect 16322 18510 16334 18562
rect 7198 18498 7250 18510
rect 8990 18498 9042 18510
rect 16718 18498 16770 18510
rect 17614 18562 17666 18574
rect 29486 18562 29538 18574
rect 37550 18562 37602 18574
rect 44046 18562 44098 18574
rect 18610 18510 18622 18562
rect 18674 18510 18686 18562
rect 30482 18510 30494 18562
rect 30546 18510 30558 18562
rect 43810 18510 43822 18562
rect 43874 18510 43886 18562
rect 49746 18510 49758 18562
rect 49810 18510 49822 18562
rect 17614 18498 17666 18510
rect 29486 18498 29538 18510
rect 37550 18498 37602 18510
rect 44046 18498 44098 18510
rect 6078 18450 6130 18462
rect 6078 18386 6130 18398
rect 6862 18450 6914 18462
rect 6862 18386 6914 18398
rect 7534 18450 7586 18462
rect 22430 18450 22482 18462
rect 27134 18450 27186 18462
rect 29374 18450 29426 18462
rect 37214 18450 37266 18462
rect 7858 18398 7870 18450
rect 7922 18398 7934 18450
rect 10434 18398 10446 18450
rect 10498 18398 10510 18450
rect 13346 18398 13358 18450
rect 13410 18398 13422 18450
rect 13682 18398 13694 18450
rect 13746 18398 13758 18450
rect 14578 18398 14590 18450
rect 14642 18398 14654 18450
rect 15474 18398 15486 18450
rect 15538 18398 15550 18450
rect 18722 18398 18734 18450
rect 18786 18398 18798 18450
rect 20066 18398 20078 18450
rect 20130 18398 20142 18450
rect 21298 18398 21310 18450
rect 21362 18398 21374 18450
rect 22642 18398 22654 18450
rect 22706 18398 22718 18450
rect 23762 18398 23774 18450
rect 23826 18398 23838 18450
rect 25442 18398 25454 18450
rect 25506 18398 25518 18450
rect 29138 18398 29150 18450
rect 29202 18398 29214 18450
rect 30370 18398 30382 18450
rect 30434 18398 30446 18450
rect 35522 18398 35534 18450
rect 35586 18398 35598 18450
rect 36530 18398 36542 18450
rect 36594 18398 36606 18450
rect 7534 18386 7586 18398
rect 22430 18386 22482 18398
rect 27134 18386 27186 18398
rect 29374 18386 29426 18398
rect 37214 18386 37266 18398
rect 37774 18450 37826 18462
rect 39230 18450 39282 18462
rect 43598 18450 43650 18462
rect 38770 18398 38782 18450
rect 38834 18398 38846 18450
rect 39442 18398 39454 18450
rect 39506 18398 39518 18450
rect 43250 18398 43262 18450
rect 43314 18398 43326 18450
rect 37774 18386 37826 18398
rect 39230 18386 39282 18398
rect 43598 18386 43650 18398
rect 45838 18450 45890 18462
rect 49634 18398 49646 18450
rect 49698 18398 49710 18450
rect 50530 18398 50542 18450
rect 50594 18398 50606 18450
rect 45838 18386 45890 18398
rect 6526 18338 6578 18350
rect 6526 18274 6578 18286
rect 9774 18338 9826 18350
rect 15262 18338 15314 18350
rect 26014 18338 26066 18350
rect 14242 18286 14254 18338
rect 14306 18286 14318 18338
rect 17714 18286 17726 18338
rect 17778 18286 17790 18338
rect 23314 18286 23326 18338
rect 23378 18286 23390 18338
rect 25554 18286 25566 18338
rect 25618 18286 25630 18338
rect 9774 18274 9826 18286
rect 15262 18274 15314 18286
rect 26014 18274 26066 18286
rect 27694 18338 27746 18350
rect 38558 18338 38610 18350
rect 28018 18286 28030 18338
rect 28082 18286 28094 18338
rect 35746 18286 35758 18338
rect 35810 18286 35822 18338
rect 37426 18286 37438 18338
rect 37490 18286 37502 18338
rect 27694 18274 27746 18286
rect 38558 18274 38610 18286
rect 40126 18338 40178 18350
rect 46846 18338 46898 18350
rect 46274 18286 46286 18338
rect 46338 18286 46350 18338
rect 40126 18274 40178 18286
rect 46846 18274 46898 18286
rect 47518 18338 47570 18350
rect 50306 18286 50318 18338
rect 50370 18286 50382 18338
rect 47518 18274 47570 18286
rect 5070 18226 5122 18238
rect 5070 18162 5122 18174
rect 17390 18226 17442 18238
rect 31166 18226 31218 18238
rect 23762 18174 23774 18226
rect 23826 18174 23838 18226
rect 29922 18174 29934 18226
rect 29986 18174 29998 18226
rect 17390 18162 17442 18174
rect 31166 18162 31218 18174
rect 31502 18226 31554 18238
rect 31502 18162 31554 18174
rect 36094 18226 36146 18238
rect 36094 18162 36146 18174
rect 36990 18226 37042 18238
rect 36990 18162 37042 18174
rect 38446 18226 38498 18238
rect 38446 18162 38498 18174
rect 47406 18226 47458 18238
rect 47406 18162 47458 18174
rect 1344 18058 58576 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 58576 18058
rect 1344 17972 58576 18006
rect 57934 17890 57986 17902
rect 9762 17838 9774 17890
rect 9826 17838 9838 17890
rect 28242 17838 28254 17890
rect 28306 17838 28318 17890
rect 34514 17838 34526 17890
rect 34578 17838 34590 17890
rect 57934 17826 57986 17838
rect 7758 17778 7810 17790
rect 23774 17778 23826 17790
rect 31502 17778 31554 17790
rect 48750 17778 48802 17790
rect 4386 17726 4398 17778
rect 4450 17726 4462 17778
rect 8642 17726 8654 17778
rect 8706 17726 8718 17778
rect 10658 17726 10670 17778
rect 10722 17775 10734 17778
rect 10994 17775 11006 17778
rect 10722 17729 11006 17775
rect 10722 17726 10734 17729
rect 10994 17726 11006 17729
rect 11058 17726 11070 17778
rect 15810 17726 15822 17778
rect 15874 17726 15886 17778
rect 24770 17726 24782 17778
rect 24834 17726 24846 17778
rect 32610 17726 32622 17778
rect 32674 17726 32686 17778
rect 34738 17726 34750 17778
rect 34802 17726 34814 17778
rect 42130 17726 42142 17778
rect 42194 17726 42206 17778
rect 45938 17726 45950 17778
rect 46002 17726 46014 17778
rect 7758 17714 7810 17726
rect 23774 17714 23826 17726
rect 31502 17714 31554 17726
rect 48750 17714 48802 17726
rect 7198 17666 7250 17678
rect 17614 17666 17666 17678
rect 5058 17614 5070 17666
rect 5122 17614 5134 17666
rect 5730 17614 5742 17666
rect 5794 17614 5806 17666
rect 8306 17614 8318 17666
rect 8370 17614 8382 17666
rect 10770 17614 10782 17666
rect 10834 17614 10846 17666
rect 11330 17614 11342 17666
rect 11394 17614 11406 17666
rect 13570 17614 13582 17666
rect 13634 17614 13646 17666
rect 14578 17614 14590 17666
rect 14642 17614 14654 17666
rect 15026 17614 15038 17666
rect 15090 17614 15102 17666
rect 7198 17602 7250 17614
rect 17614 17602 17666 17614
rect 17726 17666 17778 17678
rect 17726 17602 17778 17614
rect 17950 17666 18002 17678
rect 19070 17666 19122 17678
rect 29486 17666 29538 17678
rect 18162 17614 18174 17666
rect 18226 17614 18238 17666
rect 19282 17614 19294 17666
rect 19346 17614 19358 17666
rect 22082 17614 22094 17666
rect 22146 17614 22158 17666
rect 23090 17614 23102 17666
rect 23154 17614 23166 17666
rect 24322 17614 24334 17666
rect 24386 17614 24398 17666
rect 25890 17614 25902 17666
rect 25954 17614 25966 17666
rect 26898 17614 26910 17666
rect 26962 17614 26974 17666
rect 27234 17614 27246 17666
rect 27298 17614 27310 17666
rect 17950 17602 18002 17614
rect 19070 17602 19122 17614
rect 29486 17602 29538 17614
rect 29934 17666 29986 17678
rect 34302 17666 34354 17678
rect 30370 17614 30382 17666
rect 30434 17614 30446 17666
rect 31042 17614 31054 17666
rect 31106 17614 31118 17666
rect 32162 17614 32174 17666
rect 32226 17614 32238 17666
rect 32722 17614 32734 17666
rect 32786 17614 32798 17666
rect 29934 17602 29986 17614
rect 34302 17602 34354 17614
rect 36206 17666 36258 17678
rect 36206 17602 36258 17614
rect 41694 17666 41746 17678
rect 41694 17602 41746 17614
rect 42702 17666 42754 17678
rect 42702 17602 42754 17614
rect 43934 17666 43986 17678
rect 46510 17666 46562 17678
rect 45714 17614 45726 17666
rect 45778 17614 45790 17666
rect 43934 17602 43986 17614
rect 46510 17602 46562 17614
rect 47070 17666 47122 17678
rect 48638 17666 48690 17678
rect 51326 17666 51378 17678
rect 48066 17614 48078 17666
rect 48130 17614 48142 17666
rect 49186 17614 49198 17666
rect 49250 17614 49262 17666
rect 49522 17614 49534 17666
rect 49586 17614 49598 17666
rect 55570 17614 55582 17666
rect 55634 17614 55646 17666
rect 47070 17602 47122 17614
rect 48638 17602 48690 17614
rect 51326 17602 51378 17614
rect 1710 17554 1762 17566
rect 12910 17554 12962 17566
rect 18734 17554 18786 17566
rect 6514 17502 6526 17554
rect 6578 17502 6590 17554
rect 11218 17502 11230 17554
rect 11282 17502 11294 17554
rect 13906 17502 13918 17554
rect 13970 17502 13982 17554
rect 16818 17502 16830 17554
rect 16882 17502 16894 17554
rect 17042 17502 17054 17554
rect 17106 17502 17118 17554
rect 1710 17490 1762 17502
rect 12910 17490 12962 17502
rect 18734 17490 18786 17502
rect 21422 17554 21474 17566
rect 21422 17490 21474 17502
rect 21534 17554 21586 17566
rect 29822 17554 29874 17566
rect 35758 17554 35810 17566
rect 46846 17554 46898 17566
rect 51102 17554 51154 17566
rect 22530 17502 22542 17554
rect 22594 17502 22606 17554
rect 31714 17502 31726 17554
rect 31778 17502 31790 17554
rect 33394 17502 33406 17554
rect 33458 17502 33470 17554
rect 43026 17502 43038 17554
rect 43090 17502 43102 17554
rect 50642 17502 50654 17554
rect 50706 17502 50718 17554
rect 21534 17490 21586 17502
rect 29822 17490 29874 17502
rect 35758 17490 35810 17502
rect 46846 17490 46898 17502
rect 51102 17490 51154 17502
rect 51662 17554 51714 17566
rect 51662 17490 51714 17502
rect 21198 17442 21250 17454
rect 29710 17442 29762 17454
rect 14466 17390 14478 17442
rect 14530 17390 14542 17442
rect 20626 17390 20638 17442
rect 20690 17390 20702 17442
rect 23090 17390 23102 17442
rect 23154 17390 23166 17442
rect 21198 17378 21250 17390
rect 29710 17378 29762 17390
rect 38782 17442 38834 17454
rect 43374 17442 43426 17454
rect 51214 17442 51266 17454
rect 39106 17390 39118 17442
rect 39170 17390 39182 17442
rect 47394 17390 47406 17442
rect 47458 17390 47470 17442
rect 38782 17378 38834 17390
rect 43374 17378 43426 17390
rect 51214 17378 51266 17390
rect 1344 17274 58576 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 58576 17274
rect 1344 17188 58576 17222
rect 5182 17106 5234 17118
rect 5182 17042 5234 17054
rect 5518 17106 5570 17118
rect 5518 17042 5570 17054
rect 6078 17106 6130 17118
rect 6078 17042 6130 17054
rect 6974 17106 7026 17118
rect 6974 17042 7026 17054
rect 7758 17106 7810 17118
rect 7758 17042 7810 17054
rect 8094 17106 8146 17118
rect 8094 17042 8146 17054
rect 10110 17106 10162 17118
rect 10110 17042 10162 17054
rect 10558 17106 10610 17118
rect 10558 17042 10610 17054
rect 24782 17106 24834 17118
rect 24782 17042 24834 17054
rect 25454 17106 25506 17118
rect 25454 17042 25506 17054
rect 30942 17106 30994 17118
rect 30942 17042 30994 17054
rect 41694 17106 41746 17118
rect 41694 17042 41746 17054
rect 8654 16994 8706 17006
rect 8654 16930 8706 16942
rect 16270 16994 16322 17006
rect 18622 16994 18674 17006
rect 41470 16994 41522 17006
rect 17714 16942 17726 16994
rect 17778 16942 17790 16994
rect 17938 16942 17950 16994
rect 18002 16942 18014 16994
rect 20626 16942 20638 16994
rect 20690 16942 20702 16994
rect 23762 16942 23774 16994
rect 23826 16942 23838 16994
rect 27570 16942 27582 16994
rect 27634 16942 27646 16994
rect 29250 16942 29262 16994
rect 29314 16942 29326 16994
rect 32498 16942 32510 16994
rect 32562 16942 32574 16994
rect 37650 16942 37662 16994
rect 37714 16942 37726 16994
rect 16270 16930 16322 16942
rect 18622 16930 18674 16942
rect 41470 16930 41522 16942
rect 43822 16994 43874 17006
rect 58158 16994 58210 17006
rect 50194 16942 50206 16994
rect 50258 16942 50270 16994
rect 43822 16930 43874 16942
rect 58158 16930 58210 16942
rect 7198 16882 7250 16894
rect 11342 16882 11394 16894
rect 15486 16882 15538 16894
rect 10770 16830 10782 16882
rect 10834 16830 10846 16882
rect 14354 16830 14366 16882
rect 14418 16830 14430 16882
rect 15250 16830 15262 16882
rect 15314 16830 15326 16882
rect 7198 16818 7250 16830
rect 11342 16818 11394 16830
rect 15486 16818 15538 16830
rect 16830 16882 16882 16894
rect 16830 16818 16882 16830
rect 18510 16882 18562 16894
rect 33854 16882 33906 16894
rect 18834 16830 18846 16882
rect 18898 16830 18910 16882
rect 19506 16830 19518 16882
rect 19570 16830 19582 16882
rect 20850 16830 20862 16882
rect 20914 16830 20926 16882
rect 22754 16830 22766 16882
rect 22818 16830 22830 16882
rect 24322 16830 24334 16882
rect 24386 16830 24398 16882
rect 25778 16830 25790 16882
rect 25842 16830 25854 16882
rect 26562 16830 26574 16882
rect 26626 16830 26638 16882
rect 27122 16830 27134 16882
rect 27186 16830 27198 16882
rect 27794 16830 27806 16882
rect 27858 16830 27870 16882
rect 28690 16830 28702 16882
rect 28754 16830 28766 16882
rect 30258 16830 30270 16882
rect 30322 16830 30334 16882
rect 31826 16830 31838 16882
rect 31890 16830 31902 16882
rect 18510 16818 18562 16830
rect 33854 16818 33906 16830
rect 34078 16882 34130 16894
rect 41022 16882 41074 16894
rect 34402 16830 34414 16882
rect 34466 16830 34478 16882
rect 35410 16830 35422 16882
rect 35474 16830 35486 16882
rect 36082 16830 36094 16882
rect 36146 16830 36158 16882
rect 36418 16830 36430 16882
rect 36482 16830 36494 16882
rect 36754 16830 36766 16882
rect 36818 16830 36830 16882
rect 37538 16830 37550 16882
rect 37602 16830 37614 16882
rect 34078 16818 34130 16830
rect 41022 16818 41074 16830
rect 41806 16882 41858 16894
rect 41806 16818 41858 16830
rect 41918 16882 41970 16894
rect 43374 16882 43426 16894
rect 47182 16882 47234 16894
rect 42466 16830 42478 16882
rect 42530 16830 42542 16882
rect 45714 16830 45726 16882
rect 45778 16830 45790 16882
rect 46946 16830 46958 16882
rect 47010 16830 47022 16882
rect 51090 16830 51102 16882
rect 51154 16830 51166 16882
rect 51762 16830 51774 16882
rect 51826 16830 51838 16882
rect 53106 16830 53118 16882
rect 53170 16830 53182 16882
rect 41918 16818 41970 16830
rect 43374 16818 43426 16830
rect 47182 16818 47234 16830
rect 6526 16770 6578 16782
rect 6178 16718 6190 16770
rect 6242 16718 6254 16770
rect 5170 16606 5182 16658
rect 5234 16655 5246 16658
rect 6193 16655 6239 16718
rect 6526 16706 6578 16718
rect 11678 16770 11730 16782
rect 11678 16706 11730 16718
rect 13470 16770 13522 16782
rect 25230 16770 25282 16782
rect 14914 16718 14926 16770
rect 14978 16718 14990 16770
rect 19394 16718 19406 16770
rect 19458 16718 19470 16770
rect 25442 16718 25454 16770
rect 25506 16718 25518 16770
rect 35522 16718 35534 16770
rect 35586 16718 35598 16770
rect 37874 16718 37886 16770
rect 37938 16718 37950 16770
rect 42578 16718 42590 16770
rect 42642 16718 42654 16770
rect 45938 16718 45950 16770
rect 46002 16718 46014 16770
rect 50306 16718 50318 16770
rect 50370 16718 50382 16770
rect 13470 16706 13522 16718
rect 25230 16706 25282 16718
rect 5234 16609 6239 16655
rect 5234 16606 5246 16609
rect 14802 16606 14814 16658
rect 14866 16606 14878 16658
rect 19842 16606 19854 16658
rect 19906 16606 19918 16658
rect 26786 16606 26798 16658
rect 26850 16606 26862 16658
rect 35074 16606 35086 16658
rect 35138 16606 35150 16658
rect 46834 16606 46846 16658
rect 46898 16606 46910 16658
rect 1344 16490 58576 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 58576 16490
rect 1344 16404 58576 16438
rect 37886 16322 37938 16334
rect 57934 16322 57986 16334
rect 4274 16270 4286 16322
rect 4338 16319 4350 16322
rect 4946 16319 4958 16322
rect 4338 16273 4958 16319
rect 4338 16270 4350 16273
rect 4946 16270 4958 16273
rect 5010 16270 5022 16322
rect 10770 16270 10782 16322
rect 10834 16270 10846 16322
rect 41906 16270 41918 16322
rect 41970 16270 41982 16322
rect 37886 16258 37938 16270
rect 57934 16258 57986 16270
rect 4286 16210 4338 16222
rect 4286 16146 4338 16158
rect 5182 16210 5234 16222
rect 15262 16210 15314 16222
rect 9762 16158 9774 16210
rect 9826 16158 9838 16210
rect 10322 16158 10334 16210
rect 10386 16158 10398 16210
rect 5182 16146 5234 16158
rect 15262 16146 15314 16158
rect 16494 16210 16546 16222
rect 17154 16158 17166 16210
rect 17218 16158 17230 16210
rect 19730 16158 19742 16210
rect 19794 16158 19806 16210
rect 23426 16158 23438 16210
rect 23490 16158 23502 16210
rect 26898 16158 26910 16210
rect 26962 16158 26974 16210
rect 29698 16158 29710 16210
rect 29762 16158 29774 16210
rect 35970 16158 35982 16210
rect 36034 16158 36046 16210
rect 51202 16158 51214 16210
rect 51266 16158 51278 16210
rect 16494 16146 16546 16158
rect 7422 16098 7474 16110
rect 6962 16046 6974 16098
rect 7026 16046 7038 16098
rect 7422 16034 7474 16046
rect 7534 16098 7586 16110
rect 7534 16034 7586 16046
rect 7646 16098 7698 16110
rect 16830 16098 16882 16110
rect 20190 16098 20242 16110
rect 8866 16046 8878 16098
rect 8930 16046 8942 16098
rect 10434 16046 10446 16098
rect 10498 16046 10510 16098
rect 12338 16046 12350 16098
rect 12402 16046 12414 16098
rect 13570 16046 13582 16098
rect 13634 16046 13646 16098
rect 14466 16046 14478 16098
rect 14530 16046 14542 16098
rect 15586 16046 15598 16098
rect 15650 16046 15662 16098
rect 17826 16046 17838 16098
rect 17890 16046 17902 16098
rect 19954 16046 19966 16098
rect 20018 16046 20030 16098
rect 7646 16034 7698 16046
rect 16830 16034 16882 16046
rect 20190 16034 20242 16046
rect 20526 16098 20578 16110
rect 29262 16098 29314 16110
rect 33406 16098 33458 16110
rect 21298 16046 21310 16098
rect 21362 16046 21374 16098
rect 22418 16046 22430 16098
rect 22482 16046 22494 16098
rect 23314 16046 23326 16098
rect 23378 16046 23390 16098
rect 23986 16046 23998 16098
rect 24050 16046 24062 16098
rect 24994 16046 25006 16098
rect 25058 16046 25070 16098
rect 25890 16046 25902 16098
rect 25954 16046 25966 16098
rect 26786 16046 26798 16098
rect 26850 16046 26862 16098
rect 27794 16046 27806 16098
rect 27858 16046 27870 16098
rect 29810 16046 29822 16098
rect 29874 16046 29886 16098
rect 20526 16034 20578 16046
rect 29262 16034 29314 16046
rect 33406 16034 33458 16046
rect 33518 16098 33570 16110
rect 38670 16098 38722 16110
rect 41246 16098 41298 16110
rect 50206 16098 50258 16110
rect 34290 16046 34302 16098
rect 34354 16046 34366 16098
rect 37426 16046 37438 16098
rect 37490 16046 37502 16098
rect 39890 16046 39902 16098
rect 39954 16046 39966 16098
rect 40786 16046 40798 16098
rect 40850 16046 40862 16098
rect 41346 16046 41358 16098
rect 41410 16046 41422 16098
rect 50866 16046 50878 16098
rect 50930 16046 50942 16098
rect 55570 16046 55582 16098
rect 55634 16046 55646 16098
rect 33518 16034 33570 16046
rect 38670 16034 38722 16046
rect 41246 16034 41298 16046
rect 50206 16034 50258 16046
rect 4734 15986 4786 15998
rect 20414 15986 20466 15998
rect 27582 15986 27634 15998
rect 5842 15934 5854 15986
rect 5906 15934 5918 15986
rect 13682 15934 13694 15986
rect 13746 15934 13758 15986
rect 14578 15934 14590 15986
rect 14642 15934 14654 15986
rect 15138 15934 15150 15986
rect 15202 15934 15214 15986
rect 19842 15934 19854 15986
rect 19906 15934 19918 15986
rect 25106 15934 25118 15986
rect 25170 15934 25182 15986
rect 25778 15934 25790 15986
rect 25842 15934 25854 15986
rect 27010 15934 27022 15986
rect 27074 15934 27086 15986
rect 4734 15922 4786 15934
rect 20414 15922 20466 15934
rect 27582 15922 27634 15934
rect 33630 15986 33682 15998
rect 35758 15986 35810 15998
rect 38894 15986 38946 15998
rect 34626 15934 34638 15986
rect 34690 15934 34702 15986
rect 34850 15934 34862 15986
rect 34914 15934 34926 15986
rect 37090 15934 37102 15986
rect 37154 15934 37166 15986
rect 33630 15922 33682 15934
rect 35758 15922 35810 15934
rect 38894 15922 38946 15934
rect 39230 15986 39282 15998
rect 50094 15986 50146 15998
rect 39778 15934 39790 15986
rect 39842 15934 39854 15986
rect 42018 15934 42030 15986
rect 42082 15983 42094 15986
rect 42242 15983 42254 15986
rect 42082 15937 42254 15983
rect 42082 15934 42094 15937
rect 42242 15934 42254 15937
rect 42306 15934 42318 15986
rect 39230 15922 39282 15934
rect 50094 15922 50146 15934
rect 51550 15986 51602 15998
rect 51550 15922 51602 15934
rect 52670 15986 52722 15998
rect 52670 15922 52722 15934
rect 53006 15986 53058 15998
rect 53006 15922 53058 15934
rect 23886 15874 23938 15886
rect 8082 15822 8094 15874
rect 8146 15822 8158 15874
rect 14018 15822 14030 15874
rect 14082 15822 14094 15874
rect 23886 15810 23938 15822
rect 29374 15874 29426 15886
rect 29374 15810 29426 15822
rect 29598 15874 29650 15886
rect 29598 15810 29650 15822
rect 30270 15874 30322 15886
rect 30270 15810 30322 15822
rect 30830 15874 30882 15886
rect 30830 15810 30882 15822
rect 31166 15874 31218 15886
rect 31166 15810 31218 15822
rect 31614 15874 31666 15886
rect 31614 15810 31666 15822
rect 33182 15874 33234 15886
rect 38222 15874 38274 15886
rect 35186 15822 35198 15874
rect 35250 15822 35262 15874
rect 33182 15810 33234 15822
rect 38222 15810 38274 15822
rect 39006 15874 39058 15886
rect 39006 15810 39058 15822
rect 42366 15874 42418 15886
rect 42366 15810 42418 15822
rect 49870 15874 49922 15886
rect 49870 15810 49922 15822
rect 1344 15706 58576 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 58576 15706
rect 1344 15620 58576 15654
rect 5070 15538 5122 15550
rect 5070 15474 5122 15486
rect 5518 15538 5570 15550
rect 5518 15474 5570 15486
rect 5966 15538 6018 15550
rect 5966 15474 6018 15486
rect 9550 15538 9602 15550
rect 9550 15474 9602 15486
rect 10782 15538 10834 15550
rect 10782 15474 10834 15486
rect 11230 15538 11282 15550
rect 11230 15474 11282 15486
rect 17502 15538 17554 15550
rect 40798 15538 40850 15550
rect 28130 15486 28142 15538
rect 28194 15486 28206 15538
rect 29250 15486 29262 15538
rect 29314 15486 29326 15538
rect 30146 15486 30158 15538
rect 30210 15486 30222 15538
rect 17502 15474 17554 15486
rect 40798 15474 40850 15486
rect 41022 15538 41074 15550
rect 41022 15474 41074 15486
rect 43486 15538 43538 15550
rect 43486 15474 43538 15486
rect 45054 15538 45106 15550
rect 45054 15474 45106 15486
rect 45838 15538 45890 15550
rect 45838 15474 45890 15486
rect 46846 15538 46898 15550
rect 46846 15474 46898 15486
rect 11454 15426 11506 15438
rect 7074 15374 7086 15426
rect 7138 15374 7150 15426
rect 8418 15374 8430 15426
rect 8482 15374 8494 15426
rect 11454 15362 11506 15374
rect 12014 15426 12066 15438
rect 24670 15426 24722 15438
rect 31726 15426 31778 15438
rect 19170 15374 19182 15426
rect 19234 15374 19246 15426
rect 21410 15374 21422 15426
rect 21474 15374 21486 15426
rect 22754 15374 22766 15426
rect 22818 15374 22830 15426
rect 26898 15374 26910 15426
rect 26962 15374 26974 15426
rect 27682 15374 27694 15426
rect 27746 15374 27758 15426
rect 12014 15362 12066 15374
rect 24670 15362 24722 15374
rect 31726 15362 31778 15374
rect 35310 15426 35362 15438
rect 35310 15362 35362 15374
rect 45390 15426 45442 15438
rect 45390 15362 45442 15374
rect 46734 15426 46786 15438
rect 48302 15426 48354 15438
rect 47282 15374 47294 15426
rect 47346 15374 47358 15426
rect 47618 15374 47630 15426
rect 47682 15374 47694 15426
rect 46734 15362 46786 15374
rect 48302 15362 48354 15374
rect 50990 15426 51042 15438
rect 50990 15362 51042 15374
rect 51102 15426 51154 15438
rect 51102 15362 51154 15374
rect 53342 15426 53394 15438
rect 53342 15362 53394 15374
rect 11790 15314 11842 15326
rect 28702 15314 28754 15326
rect 7634 15262 7646 15314
rect 7698 15262 7710 15314
rect 8978 15262 8990 15314
rect 9042 15262 9054 15314
rect 12562 15262 12574 15314
rect 12626 15262 12638 15314
rect 14130 15262 14142 15314
rect 14194 15262 14206 15314
rect 15474 15262 15486 15314
rect 15538 15262 15550 15314
rect 18162 15262 18174 15314
rect 18226 15262 18238 15314
rect 18722 15262 18734 15314
rect 18786 15262 18798 15314
rect 20290 15262 20302 15314
rect 20354 15262 20366 15314
rect 21858 15262 21870 15314
rect 21922 15262 21934 15314
rect 22642 15262 22654 15314
rect 22706 15262 22718 15314
rect 23762 15262 23774 15314
rect 23826 15262 23838 15314
rect 25778 15262 25790 15314
rect 25842 15262 25854 15314
rect 26562 15262 26574 15314
rect 26626 15262 26638 15314
rect 28130 15262 28142 15314
rect 28194 15262 28206 15314
rect 11790 15250 11842 15262
rect 28702 15250 28754 15262
rect 28926 15314 28978 15326
rect 28926 15250 28978 15262
rect 29598 15314 29650 15326
rect 32958 15314 33010 15326
rect 31154 15262 31166 15314
rect 31218 15262 31230 15314
rect 31602 15262 31614 15314
rect 31666 15262 31678 15314
rect 29598 15250 29650 15262
rect 32958 15250 33010 15262
rect 33406 15314 33458 15326
rect 33406 15250 33458 15262
rect 33630 15314 33682 15326
rect 34750 15314 34802 15326
rect 37214 15314 37266 15326
rect 34402 15262 34414 15314
rect 34466 15262 34478 15314
rect 35074 15262 35086 15314
rect 35138 15262 35150 15314
rect 33630 15250 33682 15262
rect 34750 15250 34802 15262
rect 37214 15250 37266 15262
rect 37438 15314 37490 15326
rect 38110 15314 38162 15326
rect 39678 15314 39730 15326
rect 41134 15314 41186 15326
rect 37762 15262 37774 15314
rect 37826 15262 37838 15314
rect 38322 15262 38334 15314
rect 38386 15262 38398 15314
rect 38994 15262 39006 15314
rect 39058 15262 39070 15314
rect 39778 15262 39790 15314
rect 39842 15262 39854 15314
rect 37438 15250 37490 15262
rect 38110 15250 38162 15262
rect 39678 15250 39730 15262
rect 41134 15250 41186 15262
rect 42142 15314 42194 15326
rect 42142 15250 42194 15262
rect 42366 15314 42418 15326
rect 42366 15250 42418 15262
rect 42478 15314 42530 15326
rect 42478 15250 42530 15262
rect 43038 15314 43090 15326
rect 46174 15314 46226 15326
rect 51326 15314 51378 15326
rect 52670 15314 52722 15326
rect 45602 15262 45614 15314
rect 45666 15262 45678 15314
rect 46498 15262 46510 15314
rect 46562 15262 46574 15314
rect 47058 15262 47070 15314
rect 47122 15262 47134 15314
rect 51762 15262 51774 15314
rect 51826 15262 51838 15314
rect 43038 15250 43090 15262
rect 46174 15250 46226 15262
rect 51326 15250 51378 15262
rect 52670 15250 52722 15262
rect 53006 15314 53058 15326
rect 53006 15250 53058 15262
rect 6414 15202 6466 15214
rect 11902 15202 11954 15214
rect 18958 15202 19010 15214
rect 29822 15202 29874 15214
rect 9986 15150 9998 15202
rect 10050 15150 10062 15202
rect 13346 15150 13358 15202
rect 13410 15150 13422 15202
rect 15586 15150 15598 15202
rect 15650 15150 15662 15202
rect 20178 15150 20190 15202
rect 20242 15150 20254 15202
rect 22754 15150 22766 15202
rect 22818 15150 22830 15202
rect 24210 15150 24222 15202
rect 24274 15150 24286 15202
rect 25666 15150 25678 15202
rect 25730 15150 25742 15202
rect 26338 15150 26350 15202
rect 26402 15150 26414 15202
rect 6414 15138 6466 15150
rect 11902 15138 11954 15150
rect 18958 15138 19010 15150
rect 29822 15138 29874 15150
rect 30718 15202 30770 15214
rect 30718 15138 30770 15150
rect 33518 15202 33570 15214
rect 33518 15138 33570 15150
rect 33966 15202 34018 15214
rect 33966 15138 34018 15150
rect 34974 15202 35026 15214
rect 34974 15138 35026 15150
rect 41582 15202 41634 15214
rect 45826 15150 45838 15202
rect 45890 15150 45902 15202
rect 51874 15150 51886 15202
rect 51938 15150 51950 15202
rect 41582 15138 41634 15150
rect 42030 15090 42082 15102
rect 15250 15038 15262 15090
rect 15314 15038 15326 15090
rect 40226 15038 40238 15090
rect 40290 15038 40302 15090
rect 42030 15026 42082 15038
rect 1344 14922 58576 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 58576 14922
rect 1344 14836 58576 14870
rect 49870 14754 49922 14766
rect 21858 14702 21870 14754
rect 21922 14702 21934 14754
rect 33842 14702 33854 14754
rect 33906 14702 33918 14754
rect 40114 14702 40126 14754
rect 40178 14702 40190 14754
rect 49870 14690 49922 14702
rect 57934 14754 57986 14766
rect 57934 14690 57986 14702
rect 5182 14642 5234 14654
rect 5182 14578 5234 14590
rect 6638 14642 6690 14654
rect 8318 14642 8370 14654
rect 7298 14590 7310 14642
rect 7362 14590 7374 14642
rect 6638 14578 6690 14590
rect 8318 14578 8370 14590
rect 12126 14642 12178 14654
rect 28030 14642 28082 14654
rect 36318 14642 36370 14654
rect 45838 14642 45890 14654
rect 13570 14590 13582 14642
rect 13634 14590 13646 14642
rect 20626 14590 20638 14642
rect 20690 14590 20702 14642
rect 21970 14590 21982 14642
rect 22034 14590 22046 14642
rect 31490 14590 31502 14642
rect 31554 14590 31566 14642
rect 38546 14590 38558 14642
rect 38610 14590 38622 14642
rect 39778 14590 39790 14642
rect 39842 14590 39854 14642
rect 43810 14590 43822 14642
rect 43874 14590 43886 14642
rect 47058 14590 47070 14642
rect 47122 14590 47134 14642
rect 12126 14578 12178 14590
rect 28030 14578 28082 14590
rect 36318 14578 36370 14590
rect 45838 14578 45890 14590
rect 6190 14530 6242 14542
rect 17502 14530 17554 14542
rect 23550 14530 23602 14542
rect 6962 14478 6974 14530
rect 7026 14478 7038 14530
rect 7858 14478 7870 14530
rect 7922 14478 7934 14530
rect 9650 14478 9662 14530
rect 9714 14478 9726 14530
rect 10994 14478 11006 14530
rect 11058 14478 11070 14530
rect 11666 14478 11678 14530
rect 11730 14478 11742 14530
rect 12562 14478 12574 14530
rect 12626 14478 12638 14530
rect 13682 14478 13694 14530
rect 13746 14478 13758 14530
rect 15250 14478 15262 14530
rect 15314 14478 15326 14530
rect 16594 14478 16606 14530
rect 16658 14478 16670 14530
rect 18162 14478 18174 14530
rect 18226 14478 18238 14530
rect 20178 14478 20190 14530
rect 20242 14478 20254 14530
rect 21522 14478 21534 14530
rect 21586 14478 21598 14530
rect 22754 14478 22766 14530
rect 22818 14478 22830 14530
rect 6190 14466 6242 14478
rect 17502 14466 17554 14478
rect 23550 14466 23602 14478
rect 23998 14530 24050 14542
rect 23998 14466 24050 14478
rect 24334 14530 24386 14542
rect 24334 14466 24386 14478
rect 25006 14530 25058 14542
rect 35086 14530 35138 14542
rect 41134 14530 41186 14542
rect 25218 14478 25230 14530
rect 25282 14478 25294 14530
rect 26562 14478 26574 14530
rect 26626 14478 26638 14530
rect 28466 14478 28478 14530
rect 28530 14478 28542 14530
rect 31266 14478 31278 14530
rect 31330 14478 31342 14530
rect 33170 14478 33182 14530
rect 33234 14478 33246 14530
rect 34626 14478 34638 14530
rect 34690 14478 34702 14530
rect 35298 14478 35310 14530
rect 35362 14478 35374 14530
rect 37874 14478 37886 14530
rect 37938 14478 37950 14530
rect 38882 14478 38894 14530
rect 38946 14478 38958 14530
rect 39442 14478 39454 14530
rect 39506 14478 39518 14530
rect 25006 14466 25058 14478
rect 35086 14466 35138 14478
rect 41134 14466 41186 14478
rect 42142 14530 42194 14542
rect 42142 14466 42194 14478
rect 42366 14530 42418 14542
rect 43138 14478 43150 14530
rect 43202 14478 43214 14530
rect 44146 14478 44158 14530
rect 44210 14478 44222 14530
rect 45378 14478 45390 14530
rect 45442 14478 45454 14530
rect 48514 14478 48526 14530
rect 48578 14478 48590 14530
rect 55570 14478 55582 14530
rect 55634 14478 55646 14530
rect 42366 14466 42418 14478
rect 22990 14418 23042 14430
rect 8642 14366 8654 14418
rect 8706 14366 8718 14418
rect 10882 14366 10894 14418
rect 10946 14366 10958 14418
rect 11442 14366 11454 14418
rect 11506 14366 11518 14418
rect 12002 14366 12014 14418
rect 12066 14366 12078 14418
rect 13906 14366 13918 14418
rect 13970 14366 13982 14418
rect 18722 14366 18734 14418
rect 18786 14366 18798 14418
rect 22990 14354 23042 14366
rect 24782 14418 24834 14430
rect 24782 14354 24834 14366
rect 26238 14418 26290 14430
rect 27806 14418 27858 14430
rect 33630 14418 33682 14430
rect 41694 14418 41746 14430
rect 26898 14366 26910 14418
rect 26962 14366 26974 14418
rect 27122 14366 27134 14418
rect 27186 14366 27198 14418
rect 30482 14366 30494 14418
rect 30546 14366 30558 14418
rect 31714 14366 31726 14418
rect 31778 14366 31790 14418
rect 38658 14366 38670 14418
rect 38722 14366 38734 14418
rect 26238 14354 26290 14366
rect 27806 14354 27858 14366
rect 33630 14354 33682 14366
rect 41694 14354 41746 14366
rect 42254 14418 42306 14430
rect 45054 14418 45106 14430
rect 42802 14366 42814 14418
rect 42866 14366 42878 14418
rect 43250 14366 43262 14418
rect 43314 14366 43326 14418
rect 47506 14366 47518 14418
rect 47570 14366 47582 14418
rect 42254 14354 42306 14366
rect 45054 14354 45106 14366
rect 23326 14306 23378 14318
rect 17826 14254 17838 14306
rect 17890 14254 17902 14306
rect 23326 14242 23378 14254
rect 23438 14306 23490 14318
rect 23438 14242 23490 14254
rect 29486 14306 29538 14318
rect 29486 14242 29538 14254
rect 35758 14306 35810 14318
rect 35758 14242 35810 14254
rect 41470 14306 41522 14318
rect 41470 14242 41522 14254
rect 41806 14306 41858 14318
rect 41806 14242 41858 14254
rect 44830 14306 44882 14318
rect 44830 14242 44882 14254
rect 44942 14306 44994 14318
rect 44942 14242 44994 14254
rect 45726 14306 45778 14318
rect 45726 14242 45778 14254
rect 45950 14306 46002 14318
rect 45950 14242 46002 14254
rect 46174 14306 46226 14318
rect 46174 14242 46226 14254
rect 1344 14138 58576 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 58576 14138
rect 1344 14052 58576 14086
rect 6190 13970 6242 13982
rect 7758 13970 7810 13982
rect 7410 13918 7422 13970
rect 7474 13918 7486 13970
rect 6190 13906 6242 13918
rect 7758 13906 7810 13918
rect 8878 13970 8930 13982
rect 8878 13906 8930 13918
rect 9102 13970 9154 13982
rect 9102 13906 9154 13918
rect 16942 13970 16994 13982
rect 16942 13906 16994 13918
rect 21086 13970 21138 13982
rect 21086 13906 21138 13918
rect 21310 13970 21362 13982
rect 21310 13906 21362 13918
rect 25230 13970 25282 13982
rect 25230 13906 25282 13918
rect 25902 13970 25954 13982
rect 33294 13970 33346 13982
rect 31938 13918 31950 13970
rect 32002 13918 32014 13970
rect 25902 13906 25954 13918
rect 33294 13906 33346 13918
rect 44942 13970 44994 13982
rect 44942 13906 44994 13918
rect 45166 13970 45218 13982
rect 45166 13906 45218 13918
rect 47406 13970 47458 13982
rect 47406 13906 47458 13918
rect 47630 13970 47682 13982
rect 51762 13918 51774 13970
rect 51826 13918 51838 13970
rect 47630 13906 47682 13918
rect 8318 13858 8370 13870
rect 8318 13794 8370 13806
rect 8766 13858 8818 13870
rect 8766 13794 8818 13806
rect 10558 13858 10610 13870
rect 21534 13858 21586 13870
rect 28142 13858 28194 13870
rect 20514 13806 20526 13858
rect 20578 13806 20590 13858
rect 23090 13806 23102 13858
rect 23154 13806 23166 13858
rect 23986 13806 23998 13858
rect 24050 13806 24062 13858
rect 24434 13806 24446 13858
rect 24498 13806 24510 13858
rect 25554 13806 25566 13858
rect 25618 13806 25630 13858
rect 27122 13806 27134 13858
rect 27186 13806 27198 13858
rect 10558 13794 10610 13806
rect 21534 13794 21586 13806
rect 28142 13794 28194 13806
rect 30494 13858 30546 13870
rect 33182 13858 33234 13870
rect 31042 13806 31054 13858
rect 31106 13806 31118 13858
rect 30494 13794 30546 13806
rect 33182 13794 33234 13806
rect 33630 13858 33682 13870
rect 37774 13858 37826 13870
rect 39342 13858 39394 13870
rect 35074 13806 35086 13858
rect 35138 13806 35150 13858
rect 38434 13806 38446 13858
rect 38498 13806 38510 13858
rect 38658 13806 38670 13858
rect 38722 13806 38734 13858
rect 33630 13794 33682 13806
rect 37774 13794 37826 13806
rect 39342 13794 39394 13806
rect 43486 13858 43538 13870
rect 43486 13794 43538 13806
rect 43598 13858 43650 13870
rect 43598 13794 43650 13806
rect 44830 13858 44882 13870
rect 44830 13794 44882 13806
rect 45502 13858 45554 13870
rect 58158 13858 58210 13870
rect 46722 13806 46734 13858
rect 46786 13806 46798 13858
rect 52322 13806 52334 13858
rect 52386 13806 52398 13858
rect 45502 13794 45554 13806
rect 58158 13794 58210 13806
rect 6638 13746 6690 13758
rect 6638 13682 6690 13694
rect 6862 13746 6914 13758
rect 6862 13682 6914 13694
rect 7086 13746 7138 13758
rect 7086 13682 7138 13694
rect 10222 13746 10274 13758
rect 20974 13746 21026 13758
rect 30606 13746 30658 13758
rect 39006 13746 39058 13758
rect 47294 13746 47346 13758
rect 11330 13694 11342 13746
rect 11394 13694 11406 13746
rect 12674 13694 12686 13746
rect 12738 13694 12750 13746
rect 13122 13694 13134 13746
rect 13186 13694 13198 13746
rect 14914 13694 14926 13746
rect 14978 13694 14990 13746
rect 15474 13694 15486 13746
rect 15538 13694 15550 13746
rect 16258 13694 16270 13746
rect 16322 13694 16334 13746
rect 17602 13694 17614 13746
rect 17666 13694 17678 13746
rect 19170 13694 19182 13746
rect 19234 13694 19246 13746
rect 20402 13694 20414 13746
rect 20466 13694 20478 13746
rect 21858 13694 21870 13746
rect 21922 13694 21934 13746
rect 22978 13694 22990 13746
rect 23042 13694 23054 13746
rect 23762 13694 23774 13746
rect 23826 13694 23838 13746
rect 27010 13694 27022 13746
rect 27074 13694 27086 13746
rect 28466 13694 28478 13746
rect 28530 13694 28542 13746
rect 30258 13694 30270 13746
rect 30322 13694 30334 13746
rect 33842 13694 33854 13746
rect 33906 13694 33918 13746
rect 34962 13694 34974 13746
rect 35026 13694 35038 13746
rect 37314 13694 37326 13746
rect 37378 13694 37390 13746
rect 43250 13694 43262 13746
rect 43314 13694 43326 13746
rect 45826 13694 45838 13746
rect 45890 13694 45902 13746
rect 46386 13694 46398 13746
rect 46450 13694 46462 13746
rect 49858 13694 49870 13746
rect 49922 13694 49934 13746
rect 50306 13694 50318 13746
rect 50370 13694 50382 13746
rect 51314 13694 51326 13746
rect 51378 13694 51390 13746
rect 51650 13694 51662 13746
rect 51714 13694 51726 13746
rect 52210 13694 52222 13746
rect 52274 13694 52286 13746
rect 10222 13682 10274 13694
rect 20974 13682 21026 13694
rect 30606 13682 30658 13694
rect 39006 13682 39058 13694
rect 47294 13682 47346 13694
rect 10334 13634 10386 13646
rect 26014 13634 26066 13646
rect 31390 13634 31442 13646
rect 45390 13634 45442 13646
rect 10994 13582 11006 13634
rect 11058 13582 11070 13634
rect 18386 13582 18398 13634
rect 18450 13582 18462 13634
rect 19394 13582 19406 13634
rect 19458 13582 19470 13634
rect 22754 13582 22766 13634
rect 22818 13582 22830 13634
rect 28578 13582 28590 13634
rect 28642 13582 28654 13634
rect 34626 13582 34638 13634
rect 34690 13582 34702 13634
rect 36978 13582 36990 13634
rect 37042 13582 37054 13634
rect 46834 13582 46846 13634
rect 46898 13582 46910 13634
rect 50418 13582 50430 13634
rect 50482 13582 50494 13634
rect 10334 13570 10386 13582
rect 26014 13570 26066 13582
rect 31390 13570 31442 13582
rect 45390 13570 45442 13582
rect 16046 13522 16098 13534
rect 31614 13522 31666 13534
rect 13234 13470 13246 13522
rect 13298 13470 13310 13522
rect 20066 13470 20078 13522
rect 20130 13470 20142 13522
rect 16046 13458 16098 13470
rect 31614 13458 31666 13470
rect 1344 13354 58576 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 58576 13354
rect 1344 13268 58576 13302
rect 18958 13186 19010 13198
rect 32510 13186 32562 13198
rect 15138 13134 15150 13186
rect 15202 13134 15214 13186
rect 17826 13134 17838 13186
rect 17890 13134 17902 13186
rect 25106 13134 25118 13186
rect 25170 13134 25182 13186
rect 30818 13134 30830 13186
rect 30882 13183 30894 13186
rect 31602 13183 31614 13186
rect 30882 13137 31614 13183
rect 30882 13134 30894 13137
rect 31602 13134 31614 13137
rect 31666 13134 31678 13186
rect 18958 13122 19010 13134
rect 32510 13122 32562 13134
rect 42142 13186 42194 13198
rect 42142 13122 42194 13134
rect 49534 13186 49586 13198
rect 50754 13134 50766 13186
rect 50818 13134 50830 13186
rect 49534 13122 49586 13134
rect 6526 13074 6578 13086
rect 6526 13010 6578 13022
rect 7870 13074 7922 13086
rect 7870 13010 7922 13022
rect 8654 13074 8706 13086
rect 12910 13074 12962 13086
rect 27246 13074 27298 13086
rect 10098 13022 10110 13074
rect 10162 13022 10174 13074
rect 12114 13022 12126 13074
rect 12178 13022 12190 13074
rect 16594 13022 16606 13074
rect 16658 13022 16670 13074
rect 17602 13022 17614 13074
rect 17666 13022 17678 13074
rect 25218 13022 25230 13074
rect 25282 13022 25294 13074
rect 8654 13010 8706 13022
rect 12910 13010 12962 13022
rect 27246 13010 27298 13022
rect 28702 13074 28754 13086
rect 28702 13010 28754 13022
rect 32398 13074 32450 13086
rect 32398 13010 32450 13022
rect 43486 13074 43538 13086
rect 43486 13010 43538 13022
rect 48974 13074 49026 13086
rect 50194 13022 50206 13074
rect 50258 13022 50270 13074
rect 48974 13010 49026 13022
rect 6974 12962 7026 12974
rect 6974 12898 7026 12910
rect 8094 12962 8146 12974
rect 18846 12962 18898 12974
rect 26462 12962 26514 12974
rect 27582 12962 27634 12974
rect 8978 12910 8990 12962
rect 9042 12910 9054 12962
rect 11330 12910 11342 12962
rect 11394 12910 11406 12962
rect 11890 12910 11902 12962
rect 11954 12910 11966 12962
rect 14018 12910 14030 12962
rect 14082 12910 14094 12962
rect 16258 12910 16270 12962
rect 16322 12910 16334 12962
rect 19394 12910 19406 12962
rect 19458 12910 19470 12962
rect 21746 12910 21758 12962
rect 21810 12910 21822 12962
rect 22418 12910 22430 12962
rect 22482 12910 22494 12962
rect 23538 12910 23550 12962
rect 23602 12910 23614 12962
rect 24882 12910 24894 12962
rect 24946 12910 24958 12962
rect 26674 12910 26686 12962
rect 26738 12910 26750 12962
rect 8094 12898 8146 12910
rect 18846 12898 18898 12910
rect 26462 12898 26514 12910
rect 27582 12898 27634 12910
rect 28142 12962 28194 12974
rect 42030 12962 42082 12974
rect 29362 12910 29374 12962
rect 29426 12910 29438 12962
rect 32162 12910 32174 12962
rect 32226 12910 32238 12962
rect 28142 12898 28194 12910
rect 42030 12898 42082 12910
rect 42590 12962 42642 12974
rect 49198 12962 49250 12974
rect 42802 12910 42814 12962
rect 42866 12910 42878 12962
rect 50082 12910 50094 12962
rect 50146 12910 50158 12962
rect 42590 12898 42642 12910
rect 49198 12898 49250 12910
rect 7310 12850 7362 12862
rect 12462 12850 12514 12862
rect 36318 12850 36370 12862
rect 11218 12798 11230 12850
rect 11282 12798 11294 12850
rect 17378 12798 17390 12850
rect 17442 12798 17454 12850
rect 19730 12798 19742 12850
rect 19794 12798 19806 12850
rect 20178 12798 20190 12850
rect 20242 12798 20254 12850
rect 29474 12798 29486 12850
rect 29538 12798 29550 12850
rect 30034 12798 30046 12850
rect 30098 12798 30110 12850
rect 7310 12786 7362 12798
rect 12462 12786 12514 12798
rect 36318 12786 36370 12798
rect 36430 12850 36482 12862
rect 36430 12786 36482 12798
rect 41918 12850 41970 12862
rect 41918 12786 41970 12798
rect 13694 12738 13746 12750
rect 31054 12738 31106 12750
rect 20290 12686 20302 12738
rect 20354 12686 20366 12738
rect 30370 12686 30382 12738
rect 30434 12686 30446 12738
rect 13694 12674 13746 12686
rect 31054 12674 31106 12686
rect 31502 12738 31554 12750
rect 31502 12674 31554 12686
rect 35870 12738 35922 12750
rect 35870 12674 35922 12686
rect 36094 12738 36146 12750
rect 36094 12674 36146 12686
rect 41582 12738 41634 12750
rect 41582 12674 41634 12686
rect 58158 12738 58210 12750
rect 58158 12674 58210 12686
rect 1344 12570 58576 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 58576 12570
rect 1344 12484 58576 12518
rect 8206 12402 8258 12414
rect 8206 12338 8258 12350
rect 9998 12402 10050 12414
rect 9998 12338 10050 12350
rect 13246 12402 13298 12414
rect 16830 12402 16882 12414
rect 15474 12350 15486 12402
rect 15538 12350 15550 12402
rect 13246 12338 13298 12350
rect 16830 12338 16882 12350
rect 22542 12402 22594 12414
rect 23102 12402 23154 12414
rect 22754 12350 22766 12402
rect 22818 12350 22830 12402
rect 22542 12338 22594 12350
rect 23102 12338 23154 12350
rect 24222 12402 24274 12414
rect 24222 12338 24274 12350
rect 25454 12402 25506 12414
rect 25454 12338 25506 12350
rect 26350 12402 26402 12414
rect 26350 12338 26402 12350
rect 26686 12402 26738 12414
rect 26686 12338 26738 12350
rect 27358 12402 27410 12414
rect 27358 12338 27410 12350
rect 27806 12402 27858 12414
rect 27806 12338 27858 12350
rect 28254 12402 28306 12414
rect 28254 12338 28306 12350
rect 30830 12402 30882 12414
rect 30830 12338 30882 12350
rect 33294 12402 33346 12414
rect 33294 12338 33346 12350
rect 35198 12402 35250 12414
rect 35198 12338 35250 12350
rect 38446 12402 38498 12414
rect 38770 12350 38782 12402
rect 38834 12350 38846 12402
rect 50642 12350 50654 12402
rect 50706 12350 50718 12402
rect 38446 12338 38498 12350
rect 10222 12290 10274 12302
rect 14030 12290 14082 12302
rect 24446 12290 24498 12302
rect 11554 12238 11566 12290
rect 11618 12238 11630 12290
rect 11778 12238 11790 12290
rect 11842 12238 11854 12290
rect 17938 12238 17950 12290
rect 18002 12238 18014 12290
rect 21970 12238 21982 12290
rect 22034 12238 22046 12290
rect 10222 12226 10274 12238
rect 14030 12226 14082 12238
rect 24446 12226 24498 12238
rect 26126 12290 26178 12302
rect 26126 12226 26178 12238
rect 27694 12290 27746 12302
rect 27694 12226 27746 12238
rect 29598 12290 29650 12302
rect 29598 12226 29650 12238
rect 29710 12290 29762 12302
rect 29710 12226 29762 12238
rect 30270 12290 30322 12302
rect 30270 12226 30322 12238
rect 31054 12290 31106 12302
rect 31054 12226 31106 12238
rect 31502 12290 31554 12302
rect 47518 12290 47570 12302
rect 35858 12238 35870 12290
rect 35922 12238 35934 12290
rect 31502 12226 31554 12238
rect 47518 12226 47570 12238
rect 7310 12178 7362 12190
rect 7310 12114 7362 12126
rect 7534 12178 7586 12190
rect 7534 12114 7586 12126
rect 8766 12178 8818 12190
rect 15262 12178 15314 12190
rect 26014 12178 26066 12190
rect 11106 12126 11118 12178
rect 11170 12126 11182 12178
rect 12338 12126 12350 12178
rect 12402 12126 12414 12178
rect 13458 12126 13470 12178
rect 13522 12126 13534 12178
rect 18162 12126 18174 12178
rect 18226 12126 18238 12178
rect 19618 12126 19630 12178
rect 19682 12126 19694 12178
rect 21298 12126 21310 12178
rect 21362 12126 21374 12178
rect 8766 12114 8818 12126
rect 15262 12114 15314 12126
rect 26014 12114 26066 12126
rect 29934 12178 29986 12190
rect 29934 12114 29986 12126
rect 30494 12178 30546 12190
rect 30494 12114 30546 12126
rect 33182 12178 33234 12190
rect 33182 12114 33234 12126
rect 34750 12178 34802 12190
rect 39118 12178 39170 12190
rect 35970 12126 35982 12178
rect 36034 12126 36046 12178
rect 36866 12126 36878 12178
rect 36930 12126 36942 12178
rect 34750 12114 34802 12126
rect 39118 12114 39170 12126
rect 39678 12178 39730 12190
rect 39678 12114 39730 12126
rect 42366 12178 42418 12190
rect 44494 12178 44546 12190
rect 50094 12178 50146 12190
rect 43362 12126 43374 12178
rect 43426 12126 43438 12178
rect 46610 12126 46622 12178
rect 46674 12126 46686 12178
rect 42366 12114 42418 12126
rect 44494 12114 44546 12126
rect 50094 12114 50146 12126
rect 50318 12178 50370 12190
rect 50318 12114 50370 12126
rect 6638 12066 6690 12078
rect 6638 12002 6690 12014
rect 7086 12066 7138 12078
rect 7086 12002 7138 12014
rect 10782 12066 10834 12078
rect 10782 12002 10834 12014
rect 11902 12066 11954 12078
rect 11902 12002 11954 12014
rect 17502 12066 17554 12078
rect 17502 12002 17554 12014
rect 20414 12066 20466 12078
rect 20414 12002 20466 12014
rect 23774 12066 23826 12078
rect 23774 12002 23826 12014
rect 24334 12066 24386 12078
rect 29262 12066 29314 12078
rect 28690 12014 28702 12066
rect 28754 12014 28766 12066
rect 24334 12002 24386 12014
rect 29262 12002 29314 12014
rect 33854 12066 33906 12078
rect 41694 12066 41746 12078
rect 37202 12014 37214 12066
rect 37266 12014 37278 12066
rect 33854 12002 33906 12014
rect 41694 12002 41746 12014
rect 42590 12066 42642 12078
rect 44046 12066 44098 12078
rect 43586 12014 43598 12066
rect 43650 12014 43662 12066
rect 46722 12014 46734 12066
rect 46786 12014 46798 12066
rect 42590 12002 42642 12014
rect 44046 12002 44098 12014
rect 10446 11954 10498 11966
rect 7858 11902 7870 11954
rect 7922 11902 7934 11954
rect 10446 11890 10498 11902
rect 27806 11954 27858 11966
rect 27806 11890 27858 11902
rect 31166 11954 31218 11966
rect 31166 11890 31218 11902
rect 33294 11954 33346 11966
rect 36866 11902 36878 11954
rect 36930 11902 36942 11954
rect 42018 11902 42030 11954
rect 42082 11902 42094 11954
rect 33294 11890 33346 11902
rect 1344 11786 58576 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 58576 11786
rect 1344 11700 58576 11734
rect 22766 11618 22818 11630
rect 22766 11554 22818 11566
rect 23550 11618 23602 11630
rect 23550 11554 23602 11566
rect 24894 11618 24946 11630
rect 24894 11554 24946 11566
rect 25454 11618 25506 11630
rect 25454 11554 25506 11566
rect 46622 11618 46674 11630
rect 46622 11554 46674 11566
rect 7534 11506 7586 11518
rect 20750 11506 20802 11518
rect 25678 11506 25730 11518
rect 37438 11506 37490 11518
rect 41134 11506 41186 11518
rect 15026 11454 15038 11506
rect 15090 11454 15102 11506
rect 18386 11454 18398 11506
rect 18450 11454 18462 11506
rect 21746 11454 21758 11506
rect 21810 11454 21822 11506
rect 24322 11454 24334 11506
rect 24386 11454 24398 11506
rect 31378 11454 31390 11506
rect 31442 11454 31454 11506
rect 33730 11454 33742 11506
rect 33794 11454 33806 11506
rect 39666 11454 39678 11506
rect 39730 11454 39742 11506
rect 7534 11442 7586 11454
rect 20750 11442 20802 11454
rect 25678 11442 25730 11454
rect 37438 11442 37490 11454
rect 41134 11442 41186 11454
rect 43822 11506 43874 11518
rect 46398 11506 46450 11518
rect 45378 11454 45390 11506
rect 45442 11454 45454 11506
rect 43822 11442 43874 11454
rect 46398 11442 46450 11454
rect 46958 11506 47010 11518
rect 57934 11506 57986 11518
rect 50194 11454 50206 11506
rect 50258 11454 50270 11506
rect 46958 11442 47010 11454
rect 57934 11442 57986 11454
rect 9214 11394 9266 11406
rect 8418 11342 8430 11394
rect 8482 11342 8494 11394
rect 9214 11330 9266 11342
rect 9774 11394 9826 11406
rect 11902 11394 11954 11406
rect 18958 11394 19010 11406
rect 10546 11342 10558 11394
rect 10610 11342 10622 11394
rect 12786 11342 12798 11394
rect 12850 11342 12862 11394
rect 15250 11342 15262 11394
rect 15314 11342 15326 11394
rect 16034 11342 16046 11394
rect 16098 11342 16110 11394
rect 17042 11342 17054 11394
rect 17106 11342 17118 11394
rect 17378 11342 17390 11394
rect 17442 11342 17454 11394
rect 9774 11330 9826 11342
rect 11902 11330 11954 11342
rect 18958 11330 19010 11342
rect 19518 11394 19570 11406
rect 22990 11394 23042 11406
rect 22082 11342 22094 11394
rect 22146 11342 22158 11394
rect 22530 11342 22542 11394
rect 22594 11342 22606 11394
rect 19518 11330 19570 11342
rect 22990 11330 23042 11342
rect 23102 11394 23154 11406
rect 23102 11330 23154 11342
rect 23774 11394 23826 11406
rect 23774 11330 23826 11342
rect 23998 11394 24050 11406
rect 23998 11330 24050 11342
rect 24222 11394 24274 11406
rect 24222 11330 24274 11342
rect 25006 11394 25058 11406
rect 28590 11394 28642 11406
rect 34750 11394 34802 11406
rect 26450 11342 26462 11394
rect 26514 11342 26526 11394
rect 27346 11342 27358 11394
rect 27410 11342 27422 11394
rect 29362 11342 29374 11394
rect 29426 11342 29438 11394
rect 30146 11342 30158 11394
rect 30210 11342 30222 11394
rect 31042 11342 31054 11394
rect 31106 11342 31118 11394
rect 33282 11342 33294 11394
rect 33346 11342 33358 11394
rect 34066 11342 34078 11394
rect 34130 11342 34142 11394
rect 25006 11330 25058 11342
rect 28590 11330 28642 11342
rect 34750 11330 34802 11342
rect 35198 11394 35250 11406
rect 35198 11330 35250 11342
rect 35310 11394 35362 11406
rect 35310 11330 35362 11342
rect 36878 11394 36930 11406
rect 36878 11330 36930 11342
rect 37326 11394 37378 11406
rect 37326 11330 37378 11342
rect 37886 11394 37938 11406
rect 41806 11394 41858 11406
rect 43710 11394 43762 11406
rect 39442 11342 39454 11394
rect 39506 11342 39518 11394
rect 40338 11342 40350 11394
rect 40402 11342 40414 11394
rect 42242 11342 42254 11394
rect 42306 11342 42318 11394
rect 43362 11342 43374 11394
rect 43426 11342 43438 11394
rect 37886 11330 37938 11342
rect 41806 11330 41858 11342
rect 43710 11330 43762 11342
rect 47294 11394 47346 11406
rect 47294 11330 47346 11342
rect 47518 11394 47570 11406
rect 50306 11342 50318 11394
rect 50370 11342 50382 11394
rect 55570 11342 55582 11394
rect 55634 11342 55646 11394
rect 47518 11330 47570 11342
rect 8878 11282 8930 11294
rect 8878 11218 8930 11230
rect 12350 11282 12402 11294
rect 12350 11218 12402 11230
rect 19854 11282 19906 11294
rect 19854 11218 19906 11230
rect 19966 11282 20018 11294
rect 19966 11218 20018 11230
rect 24446 11282 24498 11294
rect 37998 11282 38050 11294
rect 43934 11282 43986 11294
rect 26114 11230 26126 11282
rect 26178 11279 26190 11282
rect 26450 11279 26462 11282
rect 26178 11233 26462 11279
rect 26178 11230 26190 11233
rect 26450 11230 26462 11233
rect 26514 11230 26526 11282
rect 27906 11230 27918 11282
rect 27970 11230 27982 11282
rect 30258 11230 30270 11282
rect 30322 11230 30334 11282
rect 30930 11230 30942 11282
rect 30994 11230 31006 11282
rect 34514 11230 34526 11282
rect 34578 11230 34590 11282
rect 39778 11230 39790 11282
rect 39842 11230 39854 11282
rect 42914 11230 42926 11282
rect 42978 11230 42990 11282
rect 24446 11218 24498 11230
rect 37998 11218 38050 11230
rect 43934 11218 43986 11230
rect 50990 11282 51042 11294
rect 50990 11218 51042 11230
rect 51326 11282 51378 11294
rect 51326 11218 51378 11230
rect 51662 11282 51714 11294
rect 51662 11218 51714 11230
rect 8094 11170 8146 11182
rect 13806 11170 13858 11182
rect 11218 11118 11230 11170
rect 11282 11118 11294 11170
rect 8094 11106 8146 11118
rect 13806 11106 13858 11118
rect 20190 11170 20242 11182
rect 20190 11106 20242 11118
rect 25790 11170 25842 11182
rect 32958 11170 33010 11182
rect 26562 11118 26574 11170
rect 26626 11118 26638 11170
rect 27570 11118 27582 11170
rect 27634 11118 27646 11170
rect 25790 11106 25842 11118
rect 32958 11106 33010 11118
rect 34974 11170 35026 11182
rect 34974 11106 35026 11118
rect 37550 11170 37602 11182
rect 37550 11106 37602 11118
rect 38222 11170 38274 11182
rect 38222 11106 38274 11118
rect 41470 11170 41522 11182
rect 41470 11106 41522 11118
rect 41694 11170 41746 11182
rect 45838 11170 45890 11182
rect 42354 11118 42366 11170
rect 42418 11118 42430 11170
rect 47842 11118 47854 11170
rect 47906 11118 47918 11170
rect 41694 11106 41746 11118
rect 45838 11106 45890 11118
rect 1344 11002 58576 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 58576 11002
rect 1344 10916 58576 10950
rect 8206 10834 8258 10846
rect 8206 10770 8258 10782
rect 8654 10834 8706 10846
rect 16382 10834 16434 10846
rect 14242 10782 14254 10834
rect 14306 10782 14318 10834
rect 8654 10770 8706 10782
rect 16382 10770 16434 10782
rect 17614 10834 17666 10846
rect 17614 10770 17666 10782
rect 17950 10834 18002 10846
rect 17950 10770 18002 10782
rect 22990 10834 23042 10846
rect 22990 10770 23042 10782
rect 23550 10834 23602 10846
rect 23550 10770 23602 10782
rect 24110 10834 24162 10846
rect 24110 10770 24162 10782
rect 24334 10834 24386 10846
rect 24334 10770 24386 10782
rect 24446 10834 24498 10846
rect 24446 10770 24498 10782
rect 28814 10834 28866 10846
rect 28814 10770 28866 10782
rect 29262 10834 29314 10846
rect 29262 10770 29314 10782
rect 30158 10834 30210 10846
rect 30158 10770 30210 10782
rect 34750 10834 34802 10846
rect 34750 10770 34802 10782
rect 36094 10834 36146 10846
rect 36094 10770 36146 10782
rect 36318 10834 36370 10846
rect 36318 10770 36370 10782
rect 9102 10722 9154 10734
rect 25790 10722 25842 10734
rect 34974 10722 35026 10734
rect 10210 10670 10222 10722
rect 10274 10670 10286 10722
rect 14018 10670 14030 10722
rect 14082 10670 14094 10722
rect 22530 10670 22542 10722
rect 22594 10670 22606 10722
rect 27122 10670 27134 10722
rect 27186 10670 27198 10722
rect 31490 10670 31502 10722
rect 31554 10670 31566 10722
rect 31826 10670 31838 10722
rect 31890 10670 31902 10722
rect 33730 10670 33742 10722
rect 33794 10670 33806 10722
rect 34178 10670 34190 10722
rect 34242 10670 34254 10722
rect 9102 10658 9154 10670
rect 25790 10658 25842 10670
rect 34974 10658 35026 10670
rect 57710 10722 57762 10734
rect 57710 10658 57762 10670
rect 16830 10610 16882 10622
rect 18958 10610 19010 10622
rect 10434 10558 10446 10610
rect 10498 10558 10510 10610
rect 11442 10558 11454 10610
rect 11506 10558 11518 10610
rect 12786 10558 12798 10610
rect 12850 10558 12862 10610
rect 13458 10558 13470 10610
rect 13522 10558 13534 10610
rect 15138 10558 15150 10610
rect 15202 10558 15214 10610
rect 15362 10558 15374 10610
rect 15426 10558 15438 10610
rect 15586 10558 15598 10610
rect 15650 10558 15662 10610
rect 18050 10558 18062 10610
rect 18114 10558 18126 10610
rect 16830 10546 16882 10558
rect 18958 10546 19010 10558
rect 19518 10610 19570 10622
rect 23774 10610 23826 10622
rect 29934 10610 29986 10622
rect 20738 10558 20750 10610
rect 20802 10558 20814 10610
rect 21074 10558 21086 10610
rect 21138 10558 21150 10610
rect 22194 10558 22206 10610
rect 22258 10558 22270 10610
rect 27010 10558 27022 10610
rect 27074 10558 27086 10610
rect 28130 10558 28142 10610
rect 28194 10558 28206 10610
rect 19518 10546 19570 10558
rect 23774 10546 23826 10558
rect 29934 10546 29986 10558
rect 30606 10610 30658 10622
rect 30606 10546 30658 10558
rect 33518 10610 33570 10622
rect 33518 10546 33570 10558
rect 35422 10610 35474 10622
rect 35422 10546 35474 10558
rect 35982 10610 36034 10622
rect 35982 10546 36034 10558
rect 37662 10610 37714 10622
rect 37662 10546 37714 10558
rect 38558 10610 38610 10622
rect 42142 10610 42194 10622
rect 43038 10610 43090 10622
rect 47630 10610 47682 10622
rect 38994 10558 39006 10610
rect 39058 10558 39070 10610
rect 42354 10558 42366 10610
rect 42418 10558 42430 10610
rect 46722 10558 46734 10610
rect 46786 10558 46798 10610
rect 38558 10546 38610 10558
rect 42142 10546 42194 10558
rect 43038 10546 43090 10558
rect 47630 10546 47682 10558
rect 48862 10610 48914 10622
rect 48962 10558 48974 10610
rect 49026 10558 49038 10610
rect 48862 10546 48914 10558
rect 19966 10498 20018 10510
rect 10546 10446 10558 10498
rect 10610 10446 10622 10498
rect 17938 10446 17950 10498
rect 18002 10446 18014 10498
rect 19966 10434 20018 10446
rect 20302 10498 20354 10510
rect 25342 10498 25394 10510
rect 21970 10446 21982 10498
rect 22034 10446 22046 10498
rect 20302 10434 20354 10446
rect 25342 10434 25394 10446
rect 26350 10498 26402 10510
rect 26350 10434 26402 10446
rect 26910 10498 26962 10510
rect 26910 10434 26962 10446
rect 30046 10498 30098 10510
rect 30046 10434 30098 10446
rect 31278 10498 31330 10510
rect 31278 10434 31330 10446
rect 34862 10498 34914 10510
rect 34862 10434 34914 10446
rect 37886 10498 37938 10510
rect 37886 10434 37938 10446
rect 39454 10498 39506 10510
rect 39454 10434 39506 10446
rect 41246 10498 41298 10510
rect 41246 10434 41298 10446
rect 41694 10498 41746 10510
rect 58158 10498 58210 10510
rect 47058 10446 47070 10498
rect 47122 10446 47134 10498
rect 41694 10434 41746 10446
rect 58158 10434 58210 10446
rect 30942 10386 30994 10398
rect 25218 10334 25230 10386
rect 25282 10383 25294 10386
rect 26338 10383 26350 10386
rect 25282 10337 26350 10383
rect 25282 10334 25294 10337
rect 26338 10334 26350 10337
rect 26402 10334 26414 10386
rect 30942 10322 30994 10334
rect 33182 10386 33234 10398
rect 50206 10386 50258 10398
rect 37314 10334 37326 10386
rect 37378 10334 37390 10386
rect 41234 10334 41246 10386
rect 41298 10383 41310 10386
rect 41682 10383 41694 10386
rect 41298 10337 41694 10383
rect 41298 10334 41310 10337
rect 41682 10334 41694 10337
rect 41746 10334 41758 10386
rect 33182 10322 33234 10334
rect 50206 10322 50258 10334
rect 1344 10218 58576 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 58576 10218
rect 1344 10132 58576 10166
rect 25454 10050 25506 10062
rect 25454 9986 25506 9998
rect 25790 10050 25842 10062
rect 25790 9986 25842 9998
rect 26462 10050 26514 10062
rect 26462 9986 26514 9998
rect 34302 10050 34354 10062
rect 34302 9986 34354 9998
rect 34638 10050 34690 10062
rect 34638 9986 34690 9998
rect 48974 10050 49026 10062
rect 48974 9986 49026 9998
rect 8542 9938 8594 9950
rect 8542 9874 8594 9886
rect 9438 9938 9490 9950
rect 19294 9938 19346 9950
rect 13570 9886 13582 9938
rect 13634 9886 13646 9938
rect 14690 9886 14702 9938
rect 14754 9886 14766 9938
rect 17042 9886 17054 9938
rect 17106 9886 17118 9938
rect 9438 9874 9490 9886
rect 19294 9874 19346 9886
rect 21758 9938 21810 9950
rect 21758 9874 21810 9886
rect 23326 9938 23378 9950
rect 23326 9874 23378 9886
rect 28478 9938 28530 9950
rect 35870 9938 35922 9950
rect 46286 9938 46338 9950
rect 29586 9886 29598 9938
rect 29650 9886 29662 9938
rect 40562 9886 40574 9938
rect 40626 9886 40638 9938
rect 47058 9886 47070 9938
rect 47122 9886 47134 9938
rect 28478 9874 28530 9886
rect 35870 9874 35922 9886
rect 46286 9874 46338 9886
rect 10334 9826 10386 9838
rect 9762 9774 9774 9826
rect 9826 9774 9838 9826
rect 10334 9762 10386 9774
rect 10894 9826 10946 9838
rect 15822 9826 15874 9838
rect 20638 9826 20690 9838
rect 21646 9826 21698 9838
rect 11666 9774 11678 9826
rect 11730 9774 11742 9826
rect 12226 9774 12238 9826
rect 12290 9774 12302 9826
rect 13682 9774 13694 9826
rect 13746 9774 13758 9826
rect 14914 9774 14926 9826
rect 14978 9774 14990 9826
rect 16818 9774 16830 9826
rect 16882 9774 16894 9826
rect 17266 9774 17278 9826
rect 17330 9774 17342 9826
rect 18162 9774 18174 9826
rect 18226 9774 18238 9826
rect 19170 9774 19182 9826
rect 19234 9774 19246 9826
rect 20178 9774 20190 9826
rect 20242 9774 20254 9826
rect 21298 9774 21310 9826
rect 21362 9774 21374 9826
rect 10894 9762 10946 9774
rect 15822 9762 15874 9774
rect 20638 9762 20690 9774
rect 21646 9762 21698 9774
rect 21870 9826 21922 9838
rect 22766 9826 22818 9838
rect 22194 9774 22206 9826
rect 22258 9774 22270 9826
rect 21870 9762 21922 9774
rect 22766 9762 22818 9774
rect 23438 9826 23490 9838
rect 24110 9826 24162 9838
rect 23762 9774 23774 9826
rect 23826 9774 23838 9826
rect 23438 9762 23490 9774
rect 24110 9762 24162 9774
rect 24446 9826 24498 9838
rect 27246 9826 27298 9838
rect 26450 9774 26462 9826
rect 26514 9774 26526 9826
rect 27010 9774 27022 9826
rect 27074 9774 27086 9826
rect 24446 9762 24498 9774
rect 27246 9762 27298 9774
rect 27470 9826 27522 9838
rect 29150 9826 29202 9838
rect 27682 9774 27694 9826
rect 27746 9774 27758 9826
rect 27470 9762 27522 9774
rect 29150 9762 29202 9774
rect 33406 9826 33458 9838
rect 33406 9762 33458 9774
rect 34078 9826 34130 9838
rect 34078 9762 34130 9774
rect 38782 9826 38834 9838
rect 38782 9762 38834 9774
rect 39118 9826 39170 9838
rect 40014 9826 40066 9838
rect 44046 9826 44098 9838
rect 39330 9774 39342 9826
rect 39394 9774 39406 9826
rect 40674 9774 40686 9826
rect 40738 9774 40750 9826
rect 39118 9762 39170 9774
rect 40014 9762 40066 9774
rect 44046 9762 44098 9774
rect 44158 9826 44210 9838
rect 45042 9774 45054 9826
rect 45106 9774 45118 9826
rect 46498 9774 46510 9826
rect 46562 9774 46574 9826
rect 47170 9774 47182 9826
rect 47234 9774 47246 9826
rect 44158 9762 44210 9774
rect 8990 9714 9042 9726
rect 14478 9714 14530 9726
rect 19630 9714 19682 9726
rect 11554 9662 11566 9714
rect 11618 9662 11630 9714
rect 16706 9662 16718 9714
rect 16770 9662 16782 9714
rect 18386 9662 18398 9714
rect 18450 9662 18462 9714
rect 18834 9662 18846 9714
rect 18898 9662 18910 9714
rect 8990 9650 9042 9662
rect 14478 9650 14530 9662
rect 19630 9650 19682 9662
rect 22542 9714 22594 9726
rect 22542 9650 22594 9662
rect 24222 9714 24274 9726
rect 24222 9650 24274 9662
rect 26126 9714 26178 9726
rect 26126 9650 26178 9662
rect 34526 9714 34578 9726
rect 34526 9650 34578 9662
rect 38446 9714 38498 9726
rect 38446 9650 38498 9662
rect 38558 9714 38610 9726
rect 38558 9650 38610 9662
rect 41358 9714 41410 9726
rect 49198 9714 49250 9726
rect 45378 9662 45390 9714
rect 45442 9662 45454 9714
rect 45826 9662 45838 9714
rect 45890 9662 45902 9714
rect 47842 9662 47854 9714
rect 47906 9662 47918 9714
rect 41358 9650 41410 9662
rect 49198 9650 49250 9662
rect 13022 9602 13074 9614
rect 19406 9602 19458 9614
rect 9986 9550 9998 9602
rect 10050 9550 10062 9602
rect 12114 9550 12126 9602
rect 12178 9550 12190 9602
rect 15474 9550 15486 9602
rect 15538 9550 15550 9602
rect 13022 9538 13074 9550
rect 19406 9538 19458 9550
rect 20526 9602 20578 9614
rect 20526 9538 20578 9550
rect 20750 9602 20802 9614
rect 20750 9538 20802 9550
rect 22654 9602 22706 9614
rect 22654 9538 22706 9550
rect 23214 9602 23266 9614
rect 23214 9538 23266 9550
rect 25118 9602 25170 9614
rect 25118 9538 25170 9550
rect 25678 9602 25730 9614
rect 25678 9538 25730 9550
rect 27358 9602 27410 9614
rect 27358 9538 27410 9550
rect 32398 9602 32450 9614
rect 32398 9538 32450 9550
rect 33518 9602 33570 9614
rect 33518 9538 33570 9550
rect 33630 9602 33682 9614
rect 33630 9538 33682 9550
rect 35758 9602 35810 9614
rect 35758 9538 35810 9550
rect 38222 9602 38274 9614
rect 38222 9538 38274 9550
rect 43822 9602 43874 9614
rect 43822 9538 43874 9550
rect 44270 9602 44322 9614
rect 44270 9538 44322 9550
rect 49086 9602 49138 9614
rect 49086 9538 49138 9550
rect 58158 9602 58210 9614
rect 58158 9538 58210 9550
rect 1344 9434 58576 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 58576 9434
rect 1344 9348 58576 9382
rect 9998 9266 10050 9278
rect 9998 9202 10050 9214
rect 10894 9266 10946 9278
rect 10894 9202 10946 9214
rect 11790 9266 11842 9278
rect 11790 9202 11842 9214
rect 14366 9266 14418 9278
rect 16270 9266 16322 9278
rect 15810 9214 15822 9266
rect 15874 9214 15886 9266
rect 14366 9202 14418 9214
rect 16270 9202 16322 9214
rect 16382 9266 16434 9278
rect 16382 9202 16434 9214
rect 18958 9266 19010 9278
rect 24110 9266 24162 9278
rect 23202 9214 23214 9266
rect 23266 9214 23278 9266
rect 18958 9202 19010 9214
rect 24110 9202 24162 9214
rect 26014 9266 26066 9278
rect 26014 9202 26066 9214
rect 26798 9266 26850 9278
rect 26798 9202 26850 9214
rect 27134 9266 27186 9278
rect 27134 9202 27186 9214
rect 27582 9266 27634 9278
rect 28254 9266 28306 9278
rect 27906 9214 27918 9266
rect 27970 9214 27982 9266
rect 27582 9202 27634 9214
rect 28254 9202 28306 9214
rect 28814 9266 28866 9278
rect 28814 9202 28866 9214
rect 36766 9266 36818 9278
rect 36766 9202 36818 9214
rect 39790 9266 39842 9278
rect 39790 9202 39842 9214
rect 40462 9266 40514 9278
rect 40462 9202 40514 9214
rect 45390 9266 45442 9278
rect 45390 9202 45442 9214
rect 51438 9266 51490 9278
rect 51438 9202 51490 9214
rect 13470 9154 13522 9166
rect 18510 9154 18562 9166
rect 24558 9154 24610 9166
rect 12114 9102 12126 9154
rect 12178 9102 12190 9154
rect 14914 9102 14926 9154
rect 14978 9102 14990 9154
rect 19394 9102 19406 9154
rect 19458 9102 19470 9154
rect 13470 9090 13522 9102
rect 18510 9090 18562 9102
rect 24558 9090 24610 9102
rect 26574 9154 26626 9166
rect 26574 9090 26626 9102
rect 29262 9154 29314 9166
rect 29262 9090 29314 9102
rect 29710 9154 29762 9166
rect 42590 9154 42642 9166
rect 50542 9154 50594 9166
rect 36082 9102 36094 9154
rect 36146 9102 36158 9154
rect 49074 9102 49086 9154
rect 49138 9102 49150 9154
rect 29710 9090 29762 9102
rect 42590 9090 42642 9102
rect 50542 9090 50594 9102
rect 50766 9154 50818 9166
rect 50766 9090 50818 9102
rect 10446 9042 10498 9054
rect 16494 9042 16546 9054
rect 12562 8990 12574 9042
rect 12626 8990 12638 9042
rect 14802 8990 14814 9042
rect 14866 8990 14878 9042
rect 15922 8990 15934 9042
rect 15986 8990 15998 9042
rect 10446 8978 10498 8990
rect 16494 8978 16546 8990
rect 16942 9042 16994 9054
rect 18174 9042 18226 9054
rect 19070 9042 19122 9054
rect 21982 9042 22034 9054
rect 24446 9042 24498 9054
rect 17938 8990 17950 9042
rect 18002 8990 18014 9042
rect 18722 8990 18734 9042
rect 18786 8990 18798 9042
rect 19282 8990 19294 9042
rect 19346 8990 19358 9042
rect 21634 8990 21646 9042
rect 21698 8990 21710 9042
rect 22754 8990 22766 9042
rect 22818 8990 22830 9042
rect 16942 8978 16994 8990
rect 18174 8978 18226 8990
rect 19070 8978 19122 8990
rect 21982 8978 22034 8990
rect 24446 8978 24498 8990
rect 24782 9042 24834 9054
rect 24782 8978 24834 8990
rect 25566 9042 25618 9054
rect 25566 8978 25618 8990
rect 25678 9042 25730 9054
rect 25678 8978 25730 8990
rect 25902 9042 25954 9054
rect 25902 8978 25954 8990
rect 26462 9042 26514 9054
rect 26462 8978 26514 8990
rect 31614 9042 31666 9054
rect 35310 9042 35362 9054
rect 39118 9042 39170 9054
rect 31938 8990 31950 9042
rect 32002 8990 32014 9042
rect 35970 8990 35982 9042
rect 36034 8990 36046 9042
rect 38658 8990 38670 9042
rect 38722 8990 38734 9042
rect 31614 8978 31666 8990
rect 35310 8978 35362 8990
rect 39118 8978 39170 8990
rect 39342 9042 39394 9054
rect 39342 8978 39394 8990
rect 39678 9042 39730 9054
rect 42254 9042 42306 9054
rect 41794 8990 41806 9042
rect 41858 8990 41870 9042
rect 39678 8978 39730 8990
rect 42254 8978 42306 8990
rect 42814 9042 42866 9054
rect 42814 8978 42866 8990
rect 43150 9042 43202 9054
rect 43150 8978 43202 8990
rect 44494 9042 44546 9054
rect 44494 8978 44546 8990
rect 44942 9042 44994 9054
rect 44942 8978 44994 8990
rect 45614 9042 45666 9054
rect 45614 8978 45666 8990
rect 45838 9042 45890 9054
rect 45838 8978 45890 8990
rect 46174 9042 46226 9054
rect 49410 8990 49422 9042
rect 49474 8990 49486 9042
rect 49970 8990 49982 9042
rect 50034 8990 50046 9042
rect 46174 8978 46226 8990
rect 11342 8930 11394 8942
rect 25790 8930 25842 8942
rect 12674 8878 12686 8930
rect 12738 8878 12750 8930
rect 13906 8878 13918 8930
rect 13970 8878 13982 8930
rect 11342 8866 11394 8878
rect 25790 8866 25842 8878
rect 32510 8930 32562 8942
rect 32510 8866 32562 8878
rect 43038 8930 43090 8942
rect 43038 8866 43090 8878
rect 46062 8930 46114 8942
rect 51326 8930 51378 8942
rect 49186 8878 49198 8930
rect 49250 8878 49262 8930
rect 46062 8866 46114 8878
rect 51326 8866 51378 8878
rect 13358 8818 13410 8830
rect 34974 8818 35026 8830
rect 17490 8766 17502 8818
rect 17554 8766 17566 8818
rect 28802 8766 28814 8818
rect 28866 8815 28878 8818
rect 29474 8815 29486 8818
rect 28866 8769 29486 8815
rect 28866 8766 28878 8769
rect 29474 8766 29486 8769
rect 29538 8766 29550 8818
rect 13358 8754 13410 8766
rect 34974 8754 35026 8766
rect 39790 8818 39842 8830
rect 39790 8754 39842 8766
rect 44718 8818 44770 8830
rect 44718 8754 44770 8766
rect 50878 8818 50930 8830
rect 50878 8754 50930 8766
rect 51214 8818 51266 8830
rect 51214 8754 51266 8766
rect 1344 8650 58576 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 58576 8650
rect 1344 8564 58576 8598
rect 25006 8482 25058 8494
rect 14802 8430 14814 8482
rect 14866 8430 14878 8482
rect 45826 8430 45838 8482
rect 45890 8430 45902 8482
rect 25006 8418 25058 8430
rect 10894 8370 10946 8382
rect 10894 8306 10946 8318
rect 11342 8370 11394 8382
rect 11342 8306 11394 8318
rect 21422 8370 21474 8382
rect 28254 8370 28306 8382
rect 57934 8370 57986 8382
rect 27906 8318 27918 8370
rect 27970 8318 27982 8370
rect 35298 8318 35310 8370
rect 35362 8318 35374 8370
rect 43138 8318 43150 8370
rect 43202 8318 43214 8370
rect 45490 8318 45502 8370
rect 45554 8318 45566 8370
rect 50530 8318 50542 8370
rect 50594 8318 50606 8370
rect 21422 8306 21474 8318
rect 28254 8306 28306 8318
rect 57934 8306 57986 8318
rect 11566 8258 11618 8270
rect 11566 8194 11618 8206
rect 13806 8258 13858 8270
rect 13806 8194 13858 8206
rect 14366 8258 14418 8270
rect 14366 8194 14418 8206
rect 14926 8258 14978 8270
rect 15934 8258 15986 8270
rect 15250 8206 15262 8258
rect 15314 8206 15326 8258
rect 14926 8194 14978 8206
rect 15934 8194 15986 8206
rect 16270 8258 16322 8270
rect 23774 8258 23826 8270
rect 16818 8206 16830 8258
rect 16882 8206 16894 8258
rect 18498 8206 18510 8258
rect 18562 8206 18574 8258
rect 20066 8206 20078 8258
rect 20130 8206 20142 8258
rect 23314 8206 23326 8258
rect 23378 8206 23390 8258
rect 16270 8194 16322 8206
rect 23774 8194 23826 8206
rect 23998 8258 24050 8270
rect 26910 8258 26962 8270
rect 24882 8206 24894 8258
rect 24946 8206 24958 8258
rect 23998 8194 24050 8206
rect 26910 8194 26962 8206
rect 29038 8258 29090 8270
rect 29038 8194 29090 8206
rect 29486 8258 29538 8270
rect 41470 8258 41522 8270
rect 42478 8258 42530 8270
rect 32050 8206 32062 8258
rect 32114 8206 32126 8258
rect 35522 8206 35534 8258
rect 35586 8206 35598 8258
rect 41906 8206 41918 8258
rect 41970 8206 41982 8258
rect 29486 8194 29538 8206
rect 41470 8194 41522 8206
rect 42478 8194 42530 8206
rect 42590 8258 42642 8270
rect 45154 8206 45166 8258
rect 45218 8206 45230 8258
rect 45378 8206 45390 8258
rect 45442 8206 45454 8258
rect 48178 8206 48190 8258
rect 48242 8206 48254 8258
rect 48514 8206 48526 8258
rect 48578 8206 48590 8258
rect 49522 8206 49534 8258
rect 49586 8206 49598 8258
rect 50866 8206 50878 8258
rect 50930 8206 50942 8258
rect 55570 8206 55582 8258
rect 55634 8206 55646 8258
rect 42590 8194 42642 8206
rect 27582 8146 27634 8158
rect 17490 8094 17502 8146
rect 17554 8094 17566 8146
rect 18834 8094 18846 8146
rect 18898 8094 18910 8146
rect 19954 8094 19966 8146
rect 20018 8094 20030 8146
rect 27582 8082 27634 8094
rect 27806 8146 27858 8158
rect 27806 8082 27858 8094
rect 28366 8146 28418 8158
rect 28366 8082 28418 8094
rect 28478 8146 28530 8158
rect 28478 8082 28530 8094
rect 29710 8146 29762 8158
rect 29710 8082 29762 8094
rect 30046 8146 30098 8158
rect 30046 8082 30098 8094
rect 30382 8146 30434 8158
rect 33070 8146 33122 8158
rect 32162 8094 32174 8146
rect 32226 8094 32238 8146
rect 32722 8094 32734 8146
rect 32786 8094 32798 8146
rect 30382 8082 30434 8094
rect 33070 8082 33122 8094
rect 36094 8146 36146 8158
rect 36094 8082 36146 8094
rect 38670 8146 38722 8158
rect 38670 8082 38722 8094
rect 42702 8146 42754 8158
rect 42702 8082 42754 8094
rect 48638 8146 48690 8158
rect 48638 8082 48690 8094
rect 51662 8146 51714 8158
rect 51662 8082 51714 8094
rect 51998 8146 52050 8158
rect 51998 8082 52050 8094
rect 12238 8034 12290 8046
rect 16046 8034 16098 8046
rect 11890 7982 11902 8034
rect 11954 7982 11966 8034
rect 12562 7982 12574 8034
rect 12626 7982 12638 8034
rect 12238 7970 12290 7982
rect 16046 7970 16098 7982
rect 25902 8034 25954 8046
rect 25902 7970 25954 7982
rect 26350 8034 26402 8046
rect 26350 7970 26402 7982
rect 27246 8034 27298 8046
rect 27246 7970 27298 7982
rect 29598 8034 29650 8046
rect 29598 7970 29650 7982
rect 30158 8034 30210 8046
rect 30158 7970 30210 7982
rect 33182 8034 33234 8046
rect 33182 7970 33234 7982
rect 33406 8034 33458 8046
rect 33406 7970 33458 7982
rect 38782 8034 38834 8046
rect 38782 7970 38834 7982
rect 39006 8034 39058 8046
rect 39006 7970 39058 7982
rect 1344 7866 58576 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 58576 7866
rect 1344 7780 58576 7814
rect 9886 7698 9938 7710
rect 16942 7698 16994 7710
rect 15362 7646 15374 7698
rect 15426 7646 15438 7698
rect 9886 7634 9938 7646
rect 16942 7634 16994 7646
rect 17838 7698 17890 7710
rect 17838 7634 17890 7646
rect 19854 7698 19906 7710
rect 19854 7634 19906 7646
rect 20078 7698 20130 7710
rect 20078 7634 20130 7646
rect 21534 7698 21586 7710
rect 21534 7634 21586 7646
rect 21870 7698 21922 7710
rect 21870 7634 21922 7646
rect 22542 7698 22594 7710
rect 22542 7634 22594 7646
rect 22990 7698 23042 7710
rect 22990 7634 23042 7646
rect 23438 7698 23490 7710
rect 23438 7634 23490 7646
rect 23886 7698 23938 7710
rect 23886 7634 23938 7646
rect 27358 7698 27410 7710
rect 27358 7634 27410 7646
rect 27806 7698 27858 7710
rect 27806 7634 27858 7646
rect 28254 7698 28306 7710
rect 28254 7634 28306 7646
rect 35534 7698 35586 7710
rect 35534 7634 35586 7646
rect 36094 7698 36146 7710
rect 36094 7634 36146 7646
rect 58158 7698 58210 7710
rect 58158 7634 58210 7646
rect 16382 7586 16434 7598
rect 12226 7534 12238 7586
rect 12290 7534 12302 7586
rect 14578 7534 14590 7586
rect 14642 7534 14654 7586
rect 16382 7522 16434 7534
rect 17614 7586 17666 7598
rect 17614 7522 17666 7534
rect 20190 7586 20242 7598
rect 32510 7586 32562 7598
rect 25330 7534 25342 7586
rect 25394 7534 25406 7586
rect 26002 7534 26014 7586
rect 26066 7534 26078 7586
rect 20190 7522 20242 7534
rect 32510 7522 32562 7534
rect 33406 7586 33458 7598
rect 33406 7522 33458 7534
rect 34414 7586 34466 7598
rect 34414 7522 34466 7534
rect 48974 7586 49026 7598
rect 48974 7522 49026 7534
rect 51326 7586 51378 7598
rect 51326 7522 51378 7534
rect 10222 7474 10274 7486
rect 10222 7410 10274 7422
rect 10670 7474 10722 7486
rect 10670 7410 10722 7422
rect 11006 7474 11058 7486
rect 15934 7474 15986 7486
rect 12002 7422 12014 7474
rect 12066 7422 12078 7474
rect 13458 7422 13470 7474
rect 13522 7422 13534 7474
rect 15474 7422 15486 7474
rect 15538 7422 15550 7474
rect 11006 7410 11058 7422
rect 15934 7410 15986 7422
rect 16046 7474 16098 7486
rect 20638 7474 20690 7486
rect 18610 7422 18622 7474
rect 18674 7422 18686 7474
rect 19282 7422 19294 7474
rect 19346 7422 19358 7474
rect 16046 7410 16098 7422
rect 20638 7410 20690 7422
rect 20862 7474 20914 7486
rect 20862 7410 20914 7422
rect 21646 7474 21698 7486
rect 21646 7410 21698 7422
rect 21982 7474 22034 7486
rect 21982 7410 22034 7422
rect 24222 7474 24274 7486
rect 24222 7410 24274 7422
rect 24558 7474 24610 7486
rect 35310 7474 35362 7486
rect 25666 7422 25678 7474
rect 25730 7422 25742 7474
rect 26226 7422 26238 7474
rect 26290 7422 26302 7474
rect 28914 7422 28926 7474
rect 28978 7422 28990 7474
rect 30034 7422 30046 7474
rect 30098 7422 30110 7474
rect 32050 7422 32062 7474
rect 32114 7422 32126 7474
rect 33954 7422 33966 7474
rect 34018 7422 34030 7474
rect 34850 7422 34862 7474
rect 34914 7422 34926 7474
rect 24558 7410 24610 7422
rect 35310 7410 35362 7422
rect 35646 7474 35698 7486
rect 43934 7474 43986 7486
rect 49310 7474 49362 7486
rect 51214 7474 51266 7486
rect 42242 7422 42254 7474
rect 42306 7422 42318 7474
rect 42802 7422 42814 7474
rect 42866 7422 42878 7474
rect 43362 7422 43374 7474
rect 43426 7422 43438 7474
rect 45490 7422 45502 7474
rect 45554 7422 45566 7474
rect 45826 7422 45838 7474
rect 45890 7422 45902 7474
rect 50866 7422 50878 7474
rect 50930 7422 50942 7474
rect 35646 7410 35698 7422
rect 43934 7410 43986 7422
rect 49310 7410 49362 7422
rect 51214 7410 51266 7422
rect 16270 7362 16322 7374
rect 18510 7362 18562 7374
rect 24670 7362 24722 7374
rect 17938 7310 17950 7362
rect 18002 7310 18014 7362
rect 19394 7310 19406 7362
rect 19458 7310 19470 7362
rect 16270 7298 16322 7310
rect 18510 7298 18562 7310
rect 24670 7298 24722 7310
rect 26014 7362 26066 7374
rect 26014 7298 26066 7310
rect 28814 7362 28866 7374
rect 31938 7310 31950 7362
rect 32002 7310 32014 7362
rect 34626 7310 34638 7362
rect 34690 7310 34702 7362
rect 42130 7310 42142 7362
rect 42194 7310 42206 7362
rect 47058 7310 47070 7362
rect 47122 7310 47134 7362
rect 49410 7310 49422 7362
rect 49474 7310 49486 7362
rect 28814 7298 28866 7310
rect 21086 7250 21138 7262
rect 24334 7250 24386 7262
rect 22418 7198 22430 7250
rect 22482 7247 22494 7250
rect 23090 7247 23102 7250
rect 22482 7201 23102 7247
rect 22482 7198 22494 7201
rect 23090 7198 23102 7201
rect 23154 7198 23166 7250
rect 21086 7186 21138 7198
rect 24334 7186 24386 7198
rect 29822 7250 29874 7262
rect 43586 7198 43598 7250
rect 43650 7198 43662 7250
rect 29822 7186 29874 7198
rect 1344 7082 58576 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 58576 7082
rect 1344 6996 58576 7030
rect 14030 6914 14082 6926
rect 14030 6850 14082 6862
rect 14702 6914 14754 6926
rect 25006 6914 25058 6926
rect 39118 6914 39170 6926
rect 18162 6862 18174 6914
rect 18226 6862 18238 6914
rect 35858 6862 35870 6914
rect 35922 6862 35934 6914
rect 14702 6850 14754 6862
rect 25006 6850 25058 6862
rect 39118 6850 39170 6862
rect 9886 6802 9938 6814
rect 9886 6738 9938 6750
rect 14478 6802 14530 6814
rect 19966 6802 20018 6814
rect 16146 6750 16158 6802
rect 16210 6750 16222 6802
rect 14478 6738 14530 6750
rect 19966 6738 20018 6750
rect 23102 6802 23154 6814
rect 23102 6738 23154 6750
rect 24894 6802 24946 6814
rect 29262 6802 29314 6814
rect 28354 6750 28366 6802
rect 28418 6750 28430 6802
rect 24894 6738 24946 6750
rect 29262 6738 29314 6750
rect 38558 6802 38610 6814
rect 48290 6750 48302 6802
rect 48354 6750 48366 6802
rect 38558 6738 38610 6750
rect 12238 6690 12290 6702
rect 11666 6638 11678 6690
rect 11730 6638 11742 6690
rect 12238 6626 12290 6638
rect 12798 6690 12850 6702
rect 12798 6626 12850 6638
rect 13806 6690 13858 6702
rect 13806 6626 13858 6638
rect 14254 6690 14306 6702
rect 15822 6690 15874 6702
rect 19294 6690 19346 6702
rect 20190 6690 20242 6702
rect 15026 6638 15038 6690
rect 15090 6638 15102 6690
rect 16594 6638 16606 6690
rect 16658 6638 16670 6690
rect 18386 6638 18398 6690
rect 18450 6638 18462 6690
rect 19618 6638 19630 6690
rect 19682 6638 19694 6690
rect 14254 6626 14306 6638
rect 15822 6626 15874 6638
rect 19294 6626 19346 6638
rect 20190 6626 20242 6638
rect 21422 6690 21474 6702
rect 21422 6626 21474 6638
rect 22654 6690 22706 6702
rect 22654 6626 22706 6638
rect 23998 6690 24050 6702
rect 31390 6690 31442 6702
rect 24658 6638 24670 6690
rect 24722 6638 24734 6690
rect 25330 6638 25342 6690
rect 25394 6638 25406 6690
rect 26786 6638 26798 6690
rect 26850 6638 26862 6690
rect 27458 6638 27470 6690
rect 27522 6638 27534 6690
rect 28466 6638 28478 6690
rect 28530 6638 28542 6690
rect 23998 6626 24050 6638
rect 31390 6626 31442 6638
rect 31614 6690 31666 6702
rect 31614 6626 31666 6638
rect 32062 6690 32114 6702
rect 36990 6690 37042 6702
rect 38670 6690 38722 6702
rect 32610 6638 32622 6690
rect 32674 6638 32686 6690
rect 33954 6638 33966 6690
rect 34018 6638 34030 6690
rect 35186 6638 35198 6690
rect 35250 6638 35262 6690
rect 38098 6638 38110 6690
rect 38162 6638 38174 6690
rect 32062 6626 32114 6638
rect 36990 6626 37042 6638
rect 38670 6626 38722 6638
rect 39006 6690 39058 6702
rect 49086 6690 49138 6702
rect 47842 6638 47854 6690
rect 47906 6638 47918 6690
rect 39006 6626 39058 6638
rect 49086 6626 49138 6638
rect 11342 6578 11394 6590
rect 11342 6514 11394 6526
rect 19854 6578 19906 6590
rect 19854 6514 19906 6526
rect 20414 6578 20466 6590
rect 20414 6514 20466 6526
rect 20750 6578 20802 6590
rect 20750 6514 20802 6526
rect 24446 6578 24498 6590
rect 26338 6526 26350 6578
rect 26402 6526 26414 6578
rect 28130 6526 28142 6578
rect 28194 6526 28206 6578
rect 35074 6526 35086 6578
rect 35138 6526 35150 6578
rect 24446 6514 24498 6526
rect 15150 6466 15202 6478
rect 11890 6414 11902 6466
rect 11954 6414 11966 6466
rect 15150 6402 15202 6414
rect 15486 6466 15538 6478
rect 15486 6402 15538 6414
rect 15710 6466 15762 6478
rect 15710 6402 15762 6414
rect 20638 6466 20690 6478
rect 20638 6402 20690 6414
rect 22094 6466 22146 6478
rect 25566 6466 25618 6478
rect 31502 6466 31554 6478
rect 38446 6466 38498 6478
rect 22306 6414 22318 6466
rect 22370 6414 22382 6466
rect 26450 6414 26462 6466
rect 26514 6414 26526 6466
rect 37314 6414 37326 6466
rect 37378 6414 37390 6466
rect 22094 6402 22146 6414
rect 25566 6402 25618 6414
rect 31502 6402 31554 6414
rect 38446 6402 38498 6414
rect 39118 6466 39170 6478
rect 39118 6402 39170 6414
rect 1344 6298 58576 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 58576 6298
rect 1344 6212 58576 6246
rect 12350 6130 12402 6142
rect 12350 6066 12402 6078
rect 12686 6130 12738 6142
rect 12686 6066 12738 6078
rect 13694 6130 13746 6142
rect 18622 6130 18674 6142
rect 14242 6078 14254 6130
rect 14306 6078 14318 6130
rect 13694 6066 13746 6078
rect 18622 6066 18674 6078
rect 18958 6130 19010 6142
rect 18958 6066 19010 6078
rect 20190 6130 20242 6142
rect 22094 6130 22146 6142
rect 21522 6078 21534 6130
rect 21586 6078 21598 6130
rect 20190 6066 20242 6078
rect 22094 6066 22146 6078
rect 23326 6130 23378 6142
rect 25342 6130 25394 6142
rect 23650 6078 23662 6130
rect 23714 6078 23726 6130
rect 23326 6066 23378 6078
rect 25342 6066 25394 6078
rect 25454 6130 25506 6142
rect 25454 6066 25506 6078
rect 26686 6130 26738 6142
rect 26686 6066 26738 6078
rect 26910 6130 26962 6142
rect 26910 6066 26962 6078
rect 29934 6130 29986 6142
rect 29934 6066 29986 6078
rect 30606 6130 30658 6142
rect 30606 6066 30658 6078
rect 39902 6130 39954 6142
rect 39902 6066 39954 6078
rect 41358 6130 41410 6142
rect 41358 6066 41410 6078
rect 42254 6130 42306 6142
rect 42254 6066 42306 6078
rect 44270 6130 44322 6142
rect 44270 6066 44322 6078
rect 17726 6018 17778 6030
rect 15250 5966 15262 6018
rect 15314 5966 15326 6018
rect 17726 5954 17778 5966
rect 19854 6018 19906 6030
rect 22654 6018 22706 6030
rect 20626 5966 20638 6018
rect 20690 5966 20702 6018
rect 19854 5954 19906 5966
rect 22654 5954 22706 5966
rect 24334 6018 24386 6030
rect 24334 5954 24386 5966
rect 24782 6018 24834 6030
rect 29822 6018 29874 6030
rect 28018 5966 28030 6018
rect 28082 5966 28094 6018
rect 24782 5954 24834 5966
rect 29822 5954 29874 5966
rect 31502 6018 31554 6030
rect 31502 5954 31554 5966
rect 31614 6018 31666 6030
rect 48750 6018 48802 6030
rect 35858 5966 35870 6018
rect 35922 5966 35934 6018
rect 37426 5966 37438 6018
rect 37490 5966 37502 6018
rect 31614 5954 31666 5966
rect 48750 5954 48802 5966
rect 48862 6018 48914 6030
rect 48862 5954 48914 5966
rect 50990 6018 51042 6030
rect 50990 5954 51042 5966
rect 17838 5906 17890 5918
rect 15474 5854 15486 5906
rect 15538 5854 15550 5906
rect 16258 5854 16270 5906
rect 16322 5854 16334 5906
rect 17838 5842 17890 5854
rect 18286 5906 18338 5918
rect 18286 5842 18338 5854
rect 18510 5906 18562 5918
rect 18510 5842 18562 5854
rect 19518 5906 19570 5918
rect 25230 5906 25282 5918
rect 20514 5854 20526 5906
rect 20578 5854 20590 5906
rect 21634 5854 21646 5906
rect 21698 5854 21710 5906
rect 22978 5854 22990 5906
rect 23042 5854 23054 5906
rect 19518 5842 19570 5854
rect 25230 5842 25282 5854
rect 25902 5906 25954 5918
rect 25902 5842 25954 5854
rect 26350 5906 26402 5918
rect 31838 5906 31890 5918
rect 38446 5906 38498 5918
rect 39678 5906 39730 5918
rect 27122 5854 27134 5906
rect 27186 5854 27198 5906
rect 28130 5854 28142 5906
rect 28194 5854 28206 5906
rect 29026 5854 29038 5906
rect 29090 5854 29102 5906
rect 36194 5854 36206 5906
rect 36258 5854 36270 5906
rect 39106 5854 39118 5906
rect 39170 5854 39182 5906
rect 26350 5842 26402 5854
rect 31838 5842 31890 5854
rect 38446 5842 38498 5854
rect 39678 5842 39730 5854
rect 40798 5906 40850 5918
rect 40798 5842 40850 5854
rect 41246 5906 41298 5918
rect 41246 5842 41298 5854
rect 41470 5906 41522 5918
rect 41470 5842 41522 5854
rect 41694 5906 41746 5918
rect 41694 5842 41746 5854
rect 42142 5906 42194 5918
rect 42142 5842 42194 5854
rect 42366 5906 42418 5918
rect 42366 5842 42418 5854
rect 43150 5906 43202 5918
rect 43150 5842 43202 5854
rect 43486 5906 43538 5918
rect 44606 5906 44658 5918
rect 47630 5906 47682 5918
rect 44146 5854 44158 5906
rect 44210 5854 44222 5906
rect 46722 5854 46734 5906
rect 46786 5854 46798 5906
rect 43486 5842 43538 5854
rect 44606 5842 44658 5854
rect 47630 5842 47682 5854
rect 49422 5906 49474 5918
rect 50318 5906 50370 5918
rect 49634 5854 49646 5906
rect 49698 5854 49710 5906
rect 49422 5842 49474 5854
rect 50318 5842 50370 5854
rect 50654 5906 50706 5918
rect 50654 5842 50706 5854
rect 11902 5794 11954 5806
rect 11902 5730 11954 5742
rect 13134 5794 13186 5806
rect 14814 5794 14866 5806
rect 22766 5794 22818 5806
rect 13794 5742 13806 5794
rect 13858 5742 13870 5794
rect 16146 5742 16158 5794
rect 16210 5742 16222 5794
rect 13134 5730 13186 5742
rect 14814 5730 14866 5742
rect 22766 5730 22818 5742
rect 27022 5794 27074 5806
rect 37662 5794 37714 5806
rect 45166 5794 45218 5806
rect 47294 5794 47346 5806
rect 27794 5742 27806 5794
rect 27858 5742 27870 5794
rect 29362 5742 29374 5794
rect 29426 5742 29438 5794
rect 40002 5742 40014 5794
rect 40066 5742 40078 5794
rect 43250 5742 43262 5794
rect 43314 5742 43326 5794
rect 46386 5742 46398 5794
rect 46450 5742 46462 5794
rect 27022 5730 27074 5742
rect 37662 5730 37714 5742
rect 45166 5730 45218 5742
rect 47294 5730 47346 5742
rect 13470 5682 13522 5694
rect 13470 5618 13522 5630
rect 14590 5682 14642 5694
rect 29934 5682 29986 5694
rect 42926 5682 42978 5694
rect 16482 5630 16494 5682
rect 16546 5630 16558 5682
rect 38322 5630 38334 5682
rect 38386 5630 38398 5682
rect 14590 5618 14642 5630
rect 29934 5618 29986 5630
rect 42926 5618 42978 5630
rect 43710 5682 43762 5694
rect 43710 5618 43762 5630
rect 44382 5682 44434 5694
rect 44382 5618 44434 5630
rect 45278 5682 45330 5694
rect 45278 5618 45330 5630
rect 47854 5682 47906 5694
rect 47854 5618 47906 5630
rect 48190 5682 48242 5694
rect 48190 5618 48242 5630
rect 48862 5682 48914 5694
rect 48862 5618 48914 5630
rect 1344 5514 58576 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 58576 5514
rect 1344 5428 58576 5462
rect 14814 5346 14866 5358
rect 14814 5282 14866 5294
rect 15486 5346 15538 5358
rect 15486 5282 15538 5294
rect 19854 5346 19906 5358
rect 19854 5282 19906 5294
rect 20526 5346 20578 5358
rect 20526 5282 20578 5294
rect 34750 5346 34802 5358
rect 34750 5282 34802 5294
rect 39678 5346 39730 5358
rect 39678 5282 39730 5294
rect 39902 5346 39954 5358
rect 39902 5282 39954 5294
rect 40574 5346 40626 5358
rect 40574 5282 40626 5294
rect 40798 5346 40850 5358
rect 40798 5282 40850 5294
rect 44158 5346 44210 5358
rect 13022 5234 13074 5246
rect 13022 5170 13074 5182
rect 13694 5234 13746 5246
rect 13694 5170 13746 5182
rect 14030 5234 14082 5246
rect 14030 5170 14082 5182
rect 14590 5234 14642 5246
rect 14590 5170 14642 5182
rect 16270 5234 16322 5246
rect 16270 5170 16322 5182
rect 22430 5234 22482 5246
rect 22430 5170 22482 5182
rect 23886 5234 23938 5246
rect 23886 5170 23938 5182
rect 24334 5234 24386 5246
rect 25678 5234 25730 5246
rect 25106 5182 25118 5234
rect 25170 5182 25182 5234
rect 24334 5170 24386 5182
rect 25678 5170 25730 5182
rect 26910 5234 26962 5246
rect 26910 5170 26962 5182
rect 27694 5234 27746 5246
rect 30382 5234 30434 5246
rect 40350 5234 40402 5246
rect 41570 5238 41582 5290
rect 41634 5238 41646 5290
rect 44158 5282 44210 5294
rect 46398 5346 46450 5358
rect 46398 5282 46450 5294
rect 46734 5234 46786 5246
rect 28130 5182 28142 5234
rect 28194 5182 28206 5234
rect 32722 5182 32734 5234
rect 32786 5182 32798 5234
rect 43250 5182 43262 5234
rect 43314 5182 43326 5234
rect 48066 5182 48078 5234
rect 48130 5182 48142 5234
rect 27694 5170 27746 5182
rect 30382 5170 30434 5182
rect 40350 5170 40402 5182
rect 46734 5170 46786 5182
rect 16942 5122 16994 5134
rect 15138 5070 15150 5122
rect 15202 5070 15214 5122
rect 15474 5070 15486 5122
rect 15538 5070 15550 5122
rect 16942 5058 16994 5070
rect 17614 5122 17666 5134
rect 17614 5058 17666 5070
rect 17838 5122 17890 5134
rect 17838 5058 17890 5070
rect 17950 5122 18002 5134
rect 17950 5058 18002 5070
rect 18398 5122 18450 5134
rect 18398 5058 18450 5070
rect 18622 5122 18674 5134
rect 18622 5058 18674 5070
rect 18958 5122 19010 5134
rect 18958 5058 19010 5070
rect 19742 5122 19794 5134
rect 19742 5058 19794 5070
rect 21758 5122 21810 5134
rect 21758 5058 21810 5070
rect 21982 5122 22034 5134
rect 21982 5058 22034 5070
rect 22206 5122 22258 5134
rect 22206 5058 22258 5070
rect 22654 5122 22706 5134
rect 25454 5122 25506 5134
rect 24770 5070 24782 5122
rect 24834 5070 24846 5122
rect 22654 5058 22706 5070
rect 25454 5058 25506 5070
rect 25902 5122 25954 5134
rect 25902 5058 25954 5070
rect 26014 5122 26066 5134
rect 26014 5058 26066 5070
rect 26350 5122 26402 5134
rect 26350 5058 26402 5070
rect 27022 5122 27074 5134
rect 33966 5122 34018 5134
rect 28466 5070 28478 5122
rect 28530 5070 28542 5122
rect 29138 5070 29150 5122
rect 29202 5070 29214 5122
rect 32162 5070 32174 5122
rect 32226 5070 32238 5122
rect 32834 5070 32846 5122
rect 32898 5070 32910 5122
rect 27022 5058 27074 5070
rect 33966 5058 34018 5070
rect 34526 5122 34578 5134
rect 41246 5122 41298 5134
rect 38434 5070 38446 5122
rect 38498 5070 38510 5122
rect 38658 5070 38670 5122
rect 38722 5070 38734 5122
rect 39442 5070 39454 5122
rect 39506 5070 39518 5122
rect 34526 5058 34578 5070
rect 41246 5058 41298 5070
rect 41806 5122 41858 5134
rect 45950 5122 46002 5134
rect 43026 5070 43038 5122
rect 43090 5070 43102 5122
rect 45378 5070 45390 5122
rect 45442 5070 45454 5122
rect 41806 5058 41858 5070
rect 45950 5058 46002 5070
rect 46062 5122 46114 5134
rect 46062 5058 46114 5070
rect 47070 5122 47122 5134
rect 49534 5122 49586 5134
rect 48514 5070 48526 5122
rect 48578 5070 48590 5122
rect 49074 5070 49086 5122
rect 49138 5070 49150 5122
rect 47070 5058 47122 5070
rect 49534 5058 49586 5070
rect 50094 5122 50146 5134
rect 50094 5058 50146 5070
rect 15822 5010 15874 5022
rect 15822 4946 15874 4958
rect 16606 5010 16658 5022
rect 19518 5010 19570 5022
rect 19170 4958 19182 5010
rect 19234 4958 19246 5010
rect 16606 4946 16658 4958
rect 19518 4946 19570 4958
rect 20750 5010 20802 5022
rect 20750 4946 20802 4958
rect 21422 5010 21474 5022
rect 21422 4946 21474 4958
rect 26798 5010 26850 5022
rect 34078 5010 34130 5022
rect 29362 4958 29374 5010
rect 29426 4958 29438 5010
rect 29698 4958 29710 5010
rect 29762 4958 29774 5010
rect 31826 4958 31838 5010
rect 31890 4958 31902 5010
rect 33170 4958 33182 5010
rect 33234 4958 33246 5010
rect 26798 4946 26850 4958
rect 34078 4946 34130 4958
rect 34302 5010 34354 5022
rect 34302 4946 34354 4958
rect 35646 5010 35698 5022
rect 35646 4946 35698 4958
rect 38894 5010 38946 5022
rect 38894 4946 38946 4958
rect 40014 5010 40066 5022
rect 43710 5010 43762 5022
rect 42130 4958 42142 5010
rect 42194 4958 42206 5010
rect 40014 4946 40066 4958
rect 43710 4946 43762 4958
rect 44046 5010 44098 5022
rect 44046 4946 44098 4958
rect 46510 5010 46562 5022
rect 50430 5010 50482 5022
rect 48402 4958 48414 5010
rect 48466 4958 48478 5010
rect 46510 4946 46562 4958
rect 50430 4946 50482 4958
rect 51214 5010 51266 5022
rect 51214 4946 51266 4958
rect 51326 5010 51378 5022
rect 51326 4946 51378 4958
rect 14926 4898 14978 4910
rect 14926 4834 14978 4846
rect 19070 4898 19122 4910
rect 21534 4898 21586 4910
rect 20178 4846 20190 4898
rect 20242 4846 20254 4898
rect 19070 4834 19122 4846
rect 21534 4834 21586 4846
rect 22766 4898 22818 4910
rect 22766 4834 22818 4846
rect 22878 4898 22930 4910
rect 35310 4898 35362 4910
rect 35074 4846 35086 4898
rect 35138 4846 35150 4898
rect 22878 4834 22930 4846
rect 35310 4834 35362 4846
rect 35534 4898 35586 4910
rect 35534 4834 35586 4846
rect 44158 4898 44210 4910
rect 44158 4834 44210 4846
rect 47406 4898 47458 4910
rect 47406 4834 47458 4846
rect 49422 4898 49474 4910
rect 49422 4834 49474 4846
rect 49646 4898 49698 4910
rect 49646 4834 49698 4846
rect 50766 4898 50818 4910
rect 50766 4834 50818 4846
rect 50990 4898 51042 4910
rect 50990 4834 51042 4846
rect 1344 4730 58576 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 58576 4730
rect 1344 4644 58576 4678
rect 14366 4562 14418 4574
rect 14366 4498 14418 4510
rect 15262 4562 15314 4574
rect 15262 4498 15314 4510
rect 15598 4562 15650 4574
rect 15598 4498 15650 4510
rect 16942 4562 16994 4574
rect 16942 4498 16994 4510
rect 17614 4562 17666 4574
rect 17614 4498 17666 4510
rect 18398 4562 18450 4574
rect 18398 4498 18450 4510
rect 19966 4562 20018 4574
rect 19966 4498 20018 4510
rect 21086 4562 21138 4574
rect 21086 4498 21138 4510
rect 21870 4562 21922 4574
rect 21870 4498 21922 4510
rect 23774 4562 23826 4574
rect 23774 4498 23826 4510
rect 24334 4562 24386 4574
rect 25454 4562 25506 4574
rect 24658 4510 24670 4562
rect 24722 4510 24734 4562
rect 24334 4498 24386 4510
rect 25454 4498 25506 4510
rect 26238 4562 26290 4574
rect 26238 4498 26290 4510
rect 27246 4562 27298 4574
rect 27246 4498 27298 4510
rect 28814 4562 28866 4574
rect 28814 4498 28866 4510
rect 29486 4562 29538 4574
rect 29486 4498 29538 4510
rect 30382 4562 30434 4574
rect 30382 4498 30434 4510
rect 30718 4562 30770 4574
rect 30718 4498 30770 4510
rect 30830 4562 30882 4574
rect 34078 4562 34130 4574
rect 33058 4510 33070 4562
rect 33122 4510 33134 4562
rect 30830 4498 30882 4510
rect 34078 4498 34130 4510
rect 39566 4562 39618 4574
rect 39566 4498 39618 4510
rect 42926 4562 42978 4574
rect 46834 4510 46846 4562
rect 46898 4510 46910 4562
rect 50642 4510 50654 4562
rect 50706 4510 50718 4562
rect 42926 4498 42978 4510
rect 18846 4450 18898 4462
rect 18846 4386 18898 4398
rect 19070 4450 19122 4462
rect 19070 4386 19122 4398
rect 19294 4450 19346 4462
rect 19294 4386 19346 4398
rect 22206 4450 22258 4462
rect 22206 4386 22258 4398
rect 22430 4450 22482 4462
rect 22430 4386 22482 4398
rect 23438 4450 23490 4462
rect 23438 4386 23490 4398
rect 25230 4450 25282 4462
rect 25230 4386 25282 4398
rect 28926 4450 28978 4462
rect 28926 4386 28978 4398
rect 32286 4450 32338 4462
rect 32286 4386 32338 4398
rect 33630 4450 33682 4462
rect 33630 4386 33682 4398
rect 34526 4450 34578 4462
rect 34526 4386 34578 4398
rect 39006 4450 39058 4462
rect 39006 4386 39058 4398
rect 39342 4450 39394 4462
rect 39342 4386 39394 4398
rect 42814 4450 42866 4462
rect 42814 4386 42866 4398
rect 43598 4450 43650 4462
rect 49074 4398 49086 4450
rect 49138 4398 49150 4450
rect 50754 4398 50766 4450
rect 50818 4398 50830 4450
rect 43598 4386 43650 4398
rect 19854 4338 19906 4350
rect 19854 4274 19906 4286
rect 22766 4338 22818 4350
rect 22766 4274 22818 4286
rect 30606 4338 30658 4350
rect 33406 4338 33458 4350
rect 31826 4286 31838 4338
rect 31890 4286 31902 4338
rect 30606 4274 30658 4286
rect 33406 4274 33458 4286
rect 34302 4338 34354 4350
rect 47406 4338 47458 4350
rect 35074 4286 35086 4338
rect 35138 4286 35150 4338
rect 38546 4286 38558 4338
rect 38610 4286 38622 4338
rect 43362 4286 43374 4338
rect 43426 4286 43438 4338
rect 43922 4286 43934 4338
rect 43986 4286 43998 4338
rect 51314 4286 51326 4338
rect 51378 4286 51390 4338
rect 34302 4274 34354 4286
rect 47406 4274 47458 4286
rect 14702 4226 14754 4238
rect 14702 4162 14754 4174
rect 16494 4226 16546 4238
rect 16494 4162 16546 4174
rect 19630 4226 19682 4238
rect 19630 4162 19682 4174
rect 20526 4226 20578 4238
rect 20526 4162 20578 4174
rect 21534 4226 21586 4238
rect 34414 4226 34466 4238
rect 25554 4174 25566 4226
rect 25618 4174 25630 4226
rect 31378 4174 31390 4226
rect 31442 4174 31454 4226
rect 35298 4174 35310 4226
rect 35362 4174 35374 4226
rect 38098 4174 38110 4226
rect 38162 4174 38174 4226
rect 39666 4174 39678 4226
rect 39730 4174 39742 4226
rect 48850 4174 48862 4226
rect 48914 4174 48926 4226
rect 21534 4162 21586 4174
rect 34414 4162 34466 4174
rect 22318 4114 22370 4126
rect 16482 4062 16494 4114
rect 16546 4111 16558 4114
rect 16706 4111 16718 4114
rect 16546 4065 16718 4111
rect 16546 4062 16558 4065
rect 16706 4062 16718 4065
rect 16770 4062 16782 4114
rect 22318 4050 22370 4062
rect 22990 4114 23042 4126
rect 22990 4050 23042 4062
rect 28814 4114 28866 4126
rect 44942 4114 44994 4126
rect 35858 4062 35870 4114
rect 35922 4062 35934 4114
rect 28814 4050 28866 4062
rect 44942 4050 44994 4062
rect 47182 4114 47234 4126
rect 47182 4050 47234 4062
rect 52334 4114 52386 4126
rect 52334 4050 52386 4062
rect 1344 3946 58576 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 58576 3946
rect 1344 3860 58576 3894
rect 17042 3726 17054 3778
rect 17106 3775 17118 3778
rect 18162 3775 18174 3778
rect 17106 3729 18174 3775
rect 17106 3726 17118 3729
rect 18162 3726 18174 3729
rect 18226 3726 18238 3778
rect 20738 3726 20750 3778
rect 20802 3775 20814 3778
rect 21298 3775 21310 3778
rect 20802 3729 21310 3775
rect 20802 3726 20814 3729
rect 21298 3726 21310 3729
rect 21362 3726 21374 3778
rect 14926 3666 14978 3678
rect 14926 3602 14978 3614
rect 15374 3666 15426 3678
rect 15374 3602 15426 3614
rect 15822 3666 15874 3678
rect 15822 3602 15874 3614
rect 16494 3666 16546 3678
rect 16494 3602 16546 3614
rect 17278 3666 17330 3678
rect 17278 3602 17330 3614
rect 17726 3666 17778 3678
rect 17726 3602 17778 3614
rect 18174 3666 18226 3678
rect 18174 3602 18226 3614
rect 18622 3666 18674 3678
rect 18622 3602 18674 3614
rect 19742 3666 19794 3678
rect 19742 3602 19794 3614
rect 20190 3666 20242 3678
rect 20190 3602 20242 3614
rect 20974 3666 21026 3678
rect 20974 3602 21026 3614
rect 21310 3666 21362 3678
rect 21310 3602 21362 3614
rect 22990 3666 23042 3678
rect 22990 3602 23042 3614
rect 23438 3666 23490 3678
rect 23438 3602 23490 3614
rect 28814 3666 28866 3678
rect 44606 3666 44658 3678
rect 32946 3614 32958 3666
rect 33010 3614 33022 3666
rect 28814 3602 28866 3614
rect 44606 3602 44658 3614
rect 52222 3666 52274 3678
rect 52222 3602 52274 3614
rect 19294 3554 19346 3566
rect 19294 3490 19346 3502
rect 21982 3554 22034 3566
rect 32174 3554 32226 3566
rect 38558 3554 38610 3566
rect 29026 3502 29038 3554
rect 29090 3502 29102 3554
rect 33058 3502 33070 3554
rect 33122 3502 33134 3554
rect 21982 3490 22034 3502
rect 32174 3490 32226 3502
rect 38558 3490 38610 3502
rect 38894 3554 38946 3566
rect 44034 3502 44046 3554
rect 44098 3502 44110 3554
rect 47506 3502 47518 3554
rect 47570 3502 47582 3554
rect 51426 3502 51438 3554
rect 51490 3502 51502 3554
rect 38894 3490 38946 3502
rect 38670 3442 38722 3454
rect 48962 3390 48974 3442
rect 49026 3390 49038 3442
rect 38670 3378 38722 3390
rect 5518 3330 5570 3342
rect 5518 3266 5570 3278
rect 9662 3330 9714 3342
rect 9662 3266 9714 3278
rect 30046 3330 30098 3342
rect 30046 3266 30098 3278
rect 54126 3330 54178 3342
rect 54126 3266 54178 3278
rect 1344 3162 58576 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 58576 3162
rect 1344 3076 58576 3110
<< via1 >>
rect 54462 56590 54514 56642
rect 55022 56590 55074 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 5630 56254 5682 56306
rect 6302 56254 6354 56306
rect 7646 56254 7698 56306
rect 9662 56254 9714 56306
rect 11006 56254 11058 56306
rect 11678 56254 11730 56306
rect 18286 56254 18338 56306
rect 21086 56254 21138 56306
rect 23326 56254 23378 56306
rect 27022 56254 27074 56306
rect 48414 56254 48466 56306
rect 55022 56254 55074 56306
rect 55470 56254 55522 56306
rect 13806 56142 13858 56194
rect 19182 56142 19234 56194
rect 21870 56142 21922 56194
rect 24670 56142 24722 56194
rect 25566 56142 25618 56194
rect 28478 56142 28530 56194
rect 28702 56142 28754 56194
rect 37438 56142 37490 56194
rect 19070 56030 19122 56082
rect 19742 56030 19794 56082
rect 21310 56030 21362 56082
rect 24558 56030 24610 56082
rect 30718 56030 30770 56082
rect 31502 56030 31554 56082
rect 34302 56030 34354 56082
rect 36990 56030 37042 56082
rect 42590 56030 42642 56082
rect 47406 56030 47458 56082
rect 54014 56030 54066 56082
rect 8766 55918 8818 55970
rect 14142 55918 14194 55970
rect 14702 55918 14754 55970
rect 15150 55918 15202 55970
rect 15598 55918 15650 55970
rect 16046 55918 16098 55970
rect 16494 55918 16546 55970
rect 17502 55918 17554 55970
rect 17950 55918 18002 55970
rect 18846 55918 18898 55970
rect 20078 55918 20130 55970
rect 23102 55918 23154 55970
rect 26126 55918 26178 55970
rect 26798 55918 26850 55970
rect 27582 55918 27634 55970
rect 29598 55918 29650 55970
rect 30158 55918 30210 55970
rect 31054 55918 31106 55970
rect 32398 55918 32450 55970
rect 35310 55918 35362 55970
rect 36094 55918 36146 55970
rect 36542 55918 36594 55970
rect 41022 55918 41074 55970
rect 52446 55918 52498 55970
rect 15150 55806 15202 55858
rect 16494 55806 16546 55858
rect 19182 55806 19234 55858
rect 24670 55806 24722 55858
rect 28366 55806 28418 55858
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 18062 55470 18114 55522
rect 19070 55470 19122 55522
rect 1934 55358 1986 55410
rect 14142 55358 14194 55410
rect 17838 55358 17890 55410
rect 19630 55358 19682 55410
rect 22654 55358 22706 55410
rect 24334 55358 24386 55410
rect 26798 55358 26850 55410
rect 30270 55358 30322 55410
rect 37886 55358 37938 55410
rect 47966 55358 48018 55410
rect 4174 55246 4226 55298
rect 15934 55246 15986 55298
rect 18734 55246 18786 55298
rect 19070 55246 19122 55298
rect 20750 55246 20802 55298
rect 21758 55246 21810 55298
rect 23774 55246 23826 55298
rect 23998 55246 24050 55298
rect 26686 55246 26738 55298
rect 28254 55246 28306 55298
rect 29822 55246 29874 55298
rect 31166 55246 31218 55298
rect 32174 55246 32226 55298
rect 33854 55246 33906 55298
rect 34414 55246 34466 55298
rect 35982 55246 36034 55298
rect 36206 55246 36258 55298
rect 37550 55246 37602 55298
rect 40350 55246 40402 55298
rect 40910 55246 40962 55298
rect 43374 55246 43426 55298
rect 43822 55246 43874 55298
rect 44046 55246 44098 55298
rect 44942 55246 44994 55298
rect 45278 55246 45330 55298
rect 51214 55246 51266 55298
rect 51438 55246 51490 55298
rect 15038 55134 15090 55186
rect 15374 55134 15426 55186
rect 16494 55134 16546 55186
rect 17390 55134 17442 55186
rect 22206 55134 22258 55186
rect 27918 55134 27970 55186
rect 28478 55134 28530 55186
rect 32734 55134 32786 55186
rect 33070 55134 33122 55186
rect 34862 55134 34914 55186
rect 36430 55134 36482 55186
rect 37214 55134 37266 55186
rect 38222 55134 38274 55186
rect 41022 55134 41074 55186
rect 41358 55134 41410 55186
rect 41694 55134 41746 55186
rect 42478 55134 42530 55186
rect 42702 55134 42754 55186
rect 45838 55134 45890 55186
rect 46174 55134 46226 55186
rect 46510 55134 46562 55186
rect 48190 55134 48242 55186
rect 49870 55134 49922 55186
rect 52110 55134 52162 55186
rect 52670 55134 52722 55186
rect 53006 55134 53058 55186
rect 4734 55022 4786 55074
rect 12462 55022 12514 55074
rect 12910 55022 12962 55074
rect 13918 55022 13970 55074
rect 14702 55022 14754 55074
rect 17166 55022 17218 55074
rect 17502 55022 17554 55074
rect 18398 55022 18450 55074
rect 23102 55022 23154 55074
rect 27582 55022 27634 55074
rect 28366 55022 28418 55074
rect 29262 55022 29314 55074
rect 31726 55022 31778 55074
rect 33182 55022 33234 55074
rect 33406 55022 33458 55074
rect 37326 55022 37378 55074
rect 37998 55022 38050 55074
rect 38782 55022 38834 55074
rect 39118 55022 39170 55074
rect 42254 55022 42306 55074
rect 42590 55022 42642 55074
rect 47406 55022 47458 55074
rect 50766 55022 50818 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 14926 54686 14978 54738
rect 22654 54686 22706 54738
rect 26238 54686 26290 54738
rect 45502 54686 45554 54738
rect 49982 54686 50034 54738
rect 16830 54574 16882 54626
rect 20862 54574 20914 54626
rect 21198 54574 21250 54626
rect 23662 54574 23714 54626
rect 23998 54574 24050 54626
rect 25342 54574 25394 54626
rect 33630 54574 33682 54626
rect 37662 54574 37714 54626
rect 43934 54574 43986 54626
rect 46958 54574 47010 54626
rect 49086 54574 49138 54626
rect 50766 54574 50818 54626
rect 51886 54574 51938 54626
rect 13694 54462 13746 54514
rect 14030 54462 14082 54514
rect 16606 54462 16658 54514
rect 17726 54462 17778 54514
rect 19070 54462 19122 54514
rect 19742 54462 19794 54514
rect 22430 54462 22482 54514
rect 24558 54462 24610 54514
rect 25230 54462 25282 54514
rect 26126 54462 26178 54514
rect 26910 54462 26962 54514
rect 28142 54462 28194 54514
rect 29486 54462 29538 54514
rect 30942 54462 30994 54514
rect 34526 54462 34578 54514
rect 34862 54462 34914 54514
rect 36094 54462 36146 54514
rect 36654 54462 36706 54514
rect 38222 54462 38274 54514
rect 39454 54462 39506 54514
rect 39790 54462 39842 54514
rect 41246 54462 41298 54514
rect 41806 54462 41858 54514
rect 42030 54462 42082 54514
rect 42142 54462 42194 54514
rect 42702 54462 42754 54514
rect 43374 54462 43426 54514
rect 43710 54462 43762 54514
rect 45166 54462 45218 54514
rect 46398 54462 46450 54514
rect 46846 54462 46898 54514
rect 47070 54462 47122 54514
rect 47630 54462 47682 54514
rect 48302 54462 48354 54514
rect 48750 54462 48802 54514
rect 48974 54462 49026 54514
rect 49534 54462 49586 54514
rect 50206 54462 50258 54514
rect 50654 54462 50706 54514
rect 51214 54462 51266 54514
rect 51662 54462 51714 54514
rect 53230 54462 53282 54514
rect 54574 54462 54626 54514
rect 11342 54350 11394 54402
rect 11902 54350 11954 54402
rect 12462 54350 12514 54402
rect 12910 54350 12962 54402
rect 13358 54350 13410 54402
rect 13582 54350 13634 54402
rect 14590 54350 14642 54402
rect 15486 54350 15538 54402
rect 16270 54350 16322 54402
rect 29710 54350 29762 54402
rect 31502 54350 31554 54402
rect 35422 54350 35474 54402
rect 38894 54350 38946 54402
rect 39566 54350 39618 54402
rect 41918 54350 41970 54402
rect 43822 54350 43874 54402
rect 44494 54350 44546 54402
rect 44942 54350 44994 54402
rect 47406 54350 47458 54402
rect 50990 54350 51042 54402
rect 52894 54350 52946 54402
rect 24222 54238 24274 54290
rect 31838 54238 31890 54290
rect 39006 54238 39058 54290
rect 47854 54238 47906 54290
rect 49870 54238 49922 54290
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 16382 53902 16434 53954
rect 18174 53902 18226 53954
rect 19406 53902 19458 53954
rect 34078 53902 34130 53954
rect 34302 53902 34354 53954
rect 34750 53902 34802 53954
rect 40686 53902 40738 53954
rect 41470 53902 41522 53954
rect 42814 53902 42866 53954
rect 43262 53902 43314 53954
rect 12462 53790 12514 53842
rect 18062 53790 18114 53842
rect 20414 53790 20466 53842
rect 35198 53790 35250 53842
rect 35422 53790 35474 53842
rect 40014 53790 40066 53842
rect 40798 53790 40850 53842
rect 9550 53678 9602 53730
rect 9998 53678 10050 53730
rect 12798 53678 12850 53730
rect 13918 53678 13970 53730
rect 14478 53678 14530 53730
rect 15374 53678 15426 53730
rect 15710 53678 15762 53730
rect 15934 53678 15986 53730
rect 16942 53678 16994 53730
rect 19630 53678 19682 53730
rect 20526 53678 20578 53730
rect 21534 53678 21586 53730
rect 24110 53678 24162 53730
rect 26462 53678 26514 53730
rect 26686 53678 26738 53730
rect 27694 53678 27746 53730
rect 28366 53678 28418 53730
rect 30158 53678 30210 53730
rect 30606 53678 30658 53730
rect 32286 53678 32338 53730
rect 33070 53678 33122 53730
rect 33854 53678 33906 53730
rect 35534 53678 35586 53730
rect 36878 53678 36930 53730
rect 37214 53678 37266 53730
rect 39678 53678 39730 53730
rect 42254 53678 42306 53730
rect 42478 53678 42530 53730
rect 47182 53678 47234 53730
rect 47742 53678 47794 53730
rect 47966 53678 48018 53730
rect 55582 53678 55634 53730
rect 11902 53566 11954 53618
rect 12238 53566 12290 53618
rect 17390 53566 17442 53618
rect 17838 53566 17890 53618
rect 22430 53566 22482 53618
rect 23438 53566 23490 53618
rect 28590 53566 28642 53618
rect 29150 53566 29202 53618
rect 29822 53566 29874 53618
rect 29934 53566 29986 53618
rect 31614 53566 31666 53618
rect 32174 53566 32226 53618
rect 37550 53566 37602 53618
rect 37998 53566 38050 53618
rect 40350 53566 40402 53618
rect 41358 53566 41410 53618
rect 43150 53566 43202 53618
rect 43262 53566 43314 53618
rect 47630 53566 47682 53618
rect 49086 53566 49138 53618
rect 50990 53566 51042 53618
rect 53566 53566 53618 53618
rect 53902 53566 53954 53618
rect 57262 53566 57314 53618
rect 10894 53454 10946 53506
rect 11342 53454 11394 53506
rect 13694 53454 13746 53506
rect 14814 53454 14866 53506
rect 20638 53454 20690 53506
rect 24334 53454 24386 53506
rect 27358 53454 27410 53506
rect 28030 53454 28082 53506
rect 29486 53454 29538 53506
rect 31726 53454 31778 53506
rect 33182 53454 33234 53506
rect 35982 53454 36034 53506
rect 36430 53454 36482 53506
rect 37214 53454 37266 53506
rect 39006 53454 39058 53506
rect 40910 53454 40962 53506
rect 41470 53454 41522 53506
rect 51102 53454 51154 53506
rect 51326 53454 51378 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 13358 53118 13410 53170
rect 17502 53118 17554 53170
rect 18846 53118 18898 53170
rect 22766 53118 22818 53170
rect 24334 53118 24386 53170
rect 26014 53118 26066 53170
rect 31950 53118 32002 53170
rect 32286 53118 32338 53170
rect 33630 53118 33682 53170
rect 34078 53118 34130 53170
rect 35422 53118 35474 53170
rect 37998 53118 38050 53170
rect 38894 53118 38946 53170
rect 39566 53118 39618 53170
rect 39790 53118 39842 53170
rect 40126 53118 40178 53170
rect 50878 53118 50930 53170
rect 22542 53006 22594 53058
rect 23214 53006 23266 53058
rect 23550 53006 23602 53058
rect 24670 53006 24722 53058
rect 27918 53006 27970 53058
rect 34974 53006 35026 53058
rect 39454 53006 39506 53058
rect 46510 53006 46562 53058
rect 51550 53006 51602 53058
rect 53454 53006 53506 53058
rect 10334 52894 10386 52946
rect 12126 52894 12178 52946
rect 12574 52894 12626 52946
rect 14254 52894 14306 52946
rect 15934 52894 15986 52946
rect 18510 52894 18562 52946
rect 19182 52894 19234 52946
rect 19742 52894 19794 52946
rect 21310 52894 21362 52946
rect 28478 52894 28530 52946
rect 29486 52894 29538 52946
rect 30718 52894 30770 52946
rect 45950 52894 46002 52946
rect 50094 52894 50146 52946
rect 50318 52894 50370 52946
rect 50430 52894 50482 52946
rect 52782 52894 52834 52946
rect 11454 52782 11506 52834
rect 13806 52782 13858 52834
rect 14142 52782 14194 52834
rect 16382 52782 16434 52834
rect 18062 52782 18114 52834
rect 24110 52782 24162 52834
rect 25566 52782 25618 52834
rect 26574 52782 26626 52834
rect 27022 52782 27074 52834
rect 28926 52782 28978 52834
rect 33182 52782 33234 52834
rect 34526 52782 34578 52834
rect 38446 52782 38498 52834
rect 41806 52782 41858 52834
rect 45726 52782 45778 52834
rect 51326 52782 51378 52834
rect 32958 52670 33010 52722
rect 33518 52670 33570 52722
rect 33854 52670 33906 52722
rect 34638 52670 34690 52722
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 11118 52334 11170 52386
rect 13470 52334 13522 52386
rect 13806 52334 13858 52386
rect 19406 52334 19458 52386
rect 28030 52334 28082 52386
rect 35758 52334 35810 52386
rect 41694 52334 41746 52386
rect 45838 52334 45890 52386
rect 8094 52222 8146 52274
rect 8766 52222 8818 52274
rect 9774 52222 9826 52274
rect 10670 52222 10722 52274
rect 12350 52222 12402 52274
rect 13806 52222 13858 52274
rect 17614 52222 17666 52274
rect 18286 52222 18338 52274
rect 23326 52222 23378 52274
rect 23774 52222 23826 52274
rect 27582 52222 27634 52274
rect 29598 52222 29650 52274
rect 31838 52222 31890 52274
rect 33854 52222 33906 52274
rect 37438 52222 37490 52274
rect 38558 52222 38610 52274
rect 39006 52222 39058 52274
rect 43262 52222 43314 52274
rect 44046 52222 44098 52274
rect 45278 52222 45330 52274
rect 48190 52222 48242 52274
rect 8318 52110 8370 52162
rect 9326 52110 9378 52162
rect 10446 52110 10498 52162
rect 10782 52110 10834 52162
rect 12574 52110 12626 52162
rect 14366 52110 14418 52162
rect 15822 52110 15874 52162
rect 16158 52110 16210 52162
rect 18622 52110 18674 52162
rect 20302 52110 20354 52162
rect 20414 52110 20466 52162
rect 20750 52110 20802 52162
rect 21422 52110 21474 52162
rect 22542 52110 22594 52162
rect 24222 52110 24274 52162
rect 24446 52110 24498 52162
rect 26014 52110 26066 52162
rect 27134 52110 27186 52162
rect 29038 52110 29090 52162
rect 30606 52110 30658 52162
rect 30830 52110 30882 52162
rect 31166 52110 31218 52162
rect 32174 52110 32226 52162
rect 32734 52110 32786 52162
rect 33406 52110 33458 52162
rect 34302 52110 34354 52162
rect 34526 52110 34578 52162
rect 35198 52110 35250 52162
rect 35422 52110 35474 52162
rect 37214 52110 37266 52162
rect 39454 52110 39506 52162
rect 40014 52110 40066 52162
rect 41022 52110 41074 52162
rect 41134 52110 41186 52162
rect 41246 52110 41298 52162
rect 43598 52110 43650 52162
rect 43822 52110 43874 52162
rect 44830 52110 44882 52162
rect 45726 52110 45778 52162
rect 50990 52110 51042 52162
rect 51886 52110 51938 52162
rect 12462 51998 12514 52050
rect 17166 51998 17218 52050
rect 21534 51998 21586 52050
rect 38110 51998 38162 52050
rect 40126 51998 40178 52050
rect 43486 51998 43538 52050
rect 45054 51998 45106 52050
rect 45390 51998 45442 52050
rect 51214 51998 51266 52050
rect 20638 51886 20690 51938
rect 22318 51886 22370 51938
rect 29486 51886 29538 51938
rect 29710 51886 29762 51938
rect 30382 51886 30434 51938
rect 34862 51886 34914 51938
rect 38446 51886 38498 51938
rect 39678 51886 39730 51938
rect 45838 51886 45890 51938
rect 46734 51886 46786 51938
rect 47182 51886 47234 51938
rect 47630 51886 47682 51938
rect 51998 51886 52050 51938
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 21870 51550 21922 51602
rect 22990 51550 23042 51602
rect 25230 51550 25282 51602
rect 31166 51550 31218 51602
rect 31726 51550 31778 51602
rect 39902 51550 39954 51602
rect 40126 51550 40178 51602
rect 44046 51550 44098 51602
rect 1710 51438 1762 51490
rect 9998 51438 10050 51490
rect 13918 51438 13970 51490
rect 25678 51438 25730 51490
rect 26910 51438 26962 51490
rect 29822 51438 29874 51490
rect 34862 51438 34914 51490
rect 35310 51438 35362 51490
rect 38446 51438 38498 51490
rect 39678 51438 39730 51490
rect 42702 51438 42754 51490
rect 43038 51438 43090 51490
rect 46174 51438 46226 51490
rect 50430 51438 50482 51490
rect 55022 51438 55074 51490
rect 10334 51326 10386 51378
rect 11118 51326 11170 51378
rect 12686 51326 12738 51378
rect 15486 51326 15538 51378
rect 16382 51326 16434 51378
rect 17726 51326 17778 51378
rect 18846 51326 18898 51378
rect 19182 51326 19234 51378
rect 19630 51326 19682 51378
rect 20078 51326 20130 51378
rect 20638 51326 20690 51378
rect 20750 51326 20802 51378
rect 20862 51326 20914 51378
rect 21198 51326 21250 51378
rect 21534 51326 21586 51378
rect 22542 51326 22594 51378
rect 22878 51326 22930 51378
rect 24222 51326 24274 51378
rect 25454 51326 25506 51378
rect 26126 51326 26178 51378
rect 27134 51326 27186 51378
rect 28702 51326 28754 51378
rect 29038 51326 29090 51378
rect 30718 51326 30770 51378
rect 30942 51326 30994 51378
rect 31278 51326 31330 51378
rect 33742 51326 33794 51378
rect 34190 51326 34242 51378
rect 36878 51326 36930 51378
rect 37326 51326 37378 51378
rect 40350 51326 40402 51378
rect 47518 51326 47570 51378
rect 48638 51326 48690 51378
rect 49198 51326 49250 51378
rect 49422 51326 49474 51378
rect 54686 51326 54738 51378
rect 10670 51214 10722 51266
rect 12238 51214 12290 51266
rect 13246 51214 13298 51266
rect 14254 51214 14306 51266
rect 16718 51214 16770 51266
rect 17838 51214 17890 51266
rect 23886 51214 23938 51266
rect 24558 51214 24610 51266
rect 26574 51214 26626 51266
rect 31166 51214 31218 51266
rect 32286 51214 32338 51266
rect 33182 51214 33234 51266
rect 34526 51214 34578 51266
rect 36542 51214 36594 51266
rect 43486 51214 43538 51266
rect 46510 51214 46562 51266
rect 46958 51214 47010 51266
rect 47966 51214 48018 51266
rect 14478 51102 14530 51154
rect 15598 51102 15650 51154
rect 18622 51102 18674 51154
rect 20078 51102 20130 51154
rect 22206 51102 22258 51154
rect 22542 51102 22594 51154
rect 22990 51102 23042 51154
rect 25566 51102 25618 51154
rect 32062 51102 32114 51154
rect 40238 51102 40290 51154
rect 43710 51102 43762 51154
rect 48862 51102 48914 51154
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 14142 50766 14194 50818
rect 25006 50766 25058 50818
rect 28366 50766 28418 50818
rect 29822 50766 29874 50818
rect 30158 50766 30210 50818
rect 31726 50766 31778 50818
rect 32958 50766 33010 50818
rect 37550 50766 37602 50818
rect 37998 50766 38050 50818
rect 38110 50766 38162 50818
rect 48638 50766 48690 50818
rect 52894 50766 52946 50818
rect 9550 50654 9602 50706
rect 12462 50654 12514 50706
rect 13582 50654 13634 50706
rect 15038 50654 15090 50706
rect 16718 50654 16770 50706
rect 24894 50654 24946 50706
rect 29486 50654 29538 50706
rect 30942 50654 30994 50706
rect 33294 50654 33346 50706
rect 39230 50654 39282 50706
rect 39678 50654 39730 50706
rect 43710 50654 43762 50706
rect 49646 50654 49698 50706
rect 52670 50654 52722 50706
rect 53230 50654 53282 50706
rect 53678 50654 53730 50706
rect 54574 50654 54626 50706
rect 57934 50654 57986 50706
rect 9102 50542 9154 50594
rect 13694 50542 13746 50594
rect 15598 50542 15650 50594
rect 16046 50542 16098 50594
rect 16942 50542 16994 50594
rect 17502 50542 17554 50594
rect 18398 50542 18450 50594
rect 18734 50542 18786 50594
rect 19630 50542 19682 50594
rect 20302 50542 20354 50594
rect 21310 50542 21362 50594
rect 21646 50542 21698 50594
rect 23662 50542 23714 50594
rect 24334 50542 24386 50594
rect 27358 50542 27410 50594
rect 28030 50542 28082 50594
rect 30830 50542 30882 50594
rect 31054 50542 31106 50594
rect 32286 50542 32338 50594
rect 33742 50542 33794 50594
rect 36318 50542 36370 50594
rect 37326 50542 37378 50594
rect 37998 50542 38050 50594
rect 42478 50542 42530 50594
rect 43374 50542 43426 50594
rect 45614 50542 45666 50594
rect 46174 50542 46226 50594
rect 46510 50542 46562 50594
rect 47294 50542 47346 50594
rect 48862 50542 48914 50594
rect 49086 50542 49138 50594
rect 50094 50542 50146 50594
rect 50654 50542 50706 50594
rect 53902 50542 53954 50594
rect 55582 50542 55634 50594
rect 8206 50430 8258 50482
rect 17838 50430 17890 50482
rect 19742 50430 19794 50482
rect 20750 50430 20802 50482
rect 26462 50430 26514 50482
rect 27470 50430 27522 50482
rect 30046 50430 30098 50482
rect 31390 50430 31442 50482
rect 31614 50430 31666 50482
rect 32846 50430 32898 50482
rect 35758 50430 35810 50482
rect 42142 50430 42194 50482
rect 44270 50430 44322 50482
rect 46734 50430 46786 50482
rect 46846 50430 46898 50482
rect 48078 50430 48130 50482
rect 48414 50430 48466 50482
rect 50206 50430 50258 50482
rect 50766 50430 50818 50482
rect 54910 50430 54962 50482
rect 55246 50430 55298 50482
rect 7870 50318 7922 50370
rect 8766 50318 8818 50370
rect 10334 50318 10386 50370
rect 10782 50318 10834 50370
rect 11118 50318 11170 50370
rect 11678 50318 11730 50370
rect 12014 50318 12066 50370
rect 13022 50318 13074 50370
rect 14590 50318 14642 50370
rect 18734 50318 18786 50370
rect 19966 50318 20018 50370
rect 26910 50318 26962 50370
rect 30606 50318 30658 50370
rect 32622 50318 32674 50370
rect 42814 50318 42866 50370
rect 50990 50318 51042 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 8542 49982 8594 50034
rect 15262 49982 15314 50034
rect 16830 49982 16882 50034
rect 22878 49982 22930 50034
rect 29710 49982 29762 50034
rect 31614 49982 31666 50034
rect 33630 49982 33682 50034
rect 36094 49982 36146 50034
rect 41022 49982 41074 50034
rect 41470 49982 41522 50034
rect 46958 49982 47010 50034
rect 13358 49870 13410 49922
rect 18734 49870 18786 49922
rect 20190 49870 20242 49922
rect 21422 49870 21474 49922
rect 23662 49870 23714 49922
rect 24670 49870 24722 49922
rect 26574 49870 26626 49922
rect 30382 49870 30434 49922
rect 31278 49870 31330 49922
rect 31502 49870 31554 49922
rect 32398 49870 32450 49922
rect 35198 49870 35250 49922
rect 43486 49870 43538 49922
rect 44382 49870 44434 49922
rect 46174 49870 46226 49922
rect 50990 49870 51042 49922
rect 52334 49870 52386 49922
rect 54910 49870 54962 49922
rect 8318 49758 8370 49810
rect 8878 49758 8930 49810
rect 9550 49758 9602 49810
rect 11006 49758 11058 49810
rect 11342 49758 11394 49810
rect 12350 49758 12402 49810
rect 14142 49758 14194 49810
rect 17390 49758 17442 49810
rect 17950 49758 18002 49810
rect 18510 49758 18562 49810
rect 19294 49758 19346 49810
rect 19854 49758 19906 49810
rect 21646 49758 21698 49810
rect 22766 49758 22818 49810
rect 24334 49758 24386 49810
rect 25454 49758 25506 49810
rect 27246 49758 27298 49810
rect 27806 49758 27858 49810
rect 29374 49758 29426 49810
rect 31726 49758 31778 49810
rect 31838 49758 31890 49810
rect 33518 49758 33570 49810
rect 33854 49758 33906 49810
rect 34302 49758 34354 49810
rect 35422 49758 35474 49810
rect 36654 49758 36706 49810
rect 39342 49758 39394 49810
rect 40238 49758 40290 49810
rect 42142 49758 42194 49810
rect 45278 49758 45330 49810
rect 45950 49758 46002 49810
rect 46846 49758 46898 49810
rect 51774 49758 51826 49810
rect 53902 49758 53954 49810
rect 54350 49758 54402 49810
rect 8990 49646 9042 49698
rect 9998 49646 10050 49698
rect 11454 49646 11506 49698
rect 12014 49646 12066 49698
rect 14702 49646 14754 49698
rect 15822 49646 15874 49698
rect 16382 49646 16434 49698
rect 18286 49646 18338 49698
rect 19966 49646 20018 49698
rect 34302 49646 34354 49698
rect 34974 49646 35026 49698
rect 37998 49646 38050 49698
rect 39790 49646 39842 49698
rect 50878 49646 50930 49698
rect 54014 49646 54066 49698
rect 33966 49534 34018 49586
rect 45166 49534 45218 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 9886 49198 9938 49250
rect 1934 49086 1986 49138
rect 10558 49086 10610 49138
rect 11006 49086 11058 49138
rect 16830 49086 16882 49138
rect 20190 49086 20242 49138
rect 22430 49086 22482 49138
rect 24222 49086 24274 49138
rect 26798 49086 26850 49138
rect 29486 49086 29538 49138
rect 30718 49086 30770 49138
rect 32510 49086 32562 49138
rect 32958 49086 33010 49138
rect 33518 49198 33570 49250
rect 39006 49198 39058 49250
rect 36430 49086 36482 49138
rect 37326 49086 37378 49138
rect 39790 49086 39842 49138
rect 41694 49086 41746 49138
rect 43710 49086 43762 49138
rect 44830 49086 44882 49138
rect 53118 49086 53170 49138
rect 53902 49086 53954 49138
rect 57822 49086 57874 49138
rect 4286 48974 4338 49026
rect 7422 48974 7474 49026
rect 7870 48974 7922 49026
rect 9214 48974 9266 49026
rect 9550 48974 9602 49026
rect 9774 48974 9826 49026
rect 11790 48974 11842 49026
rect 12238 48974 12290 49026
rect 12574 48974 12626 49026
rect 13022 48974 13074 49026
rect 13582 48974 13634 49026
rect 13918 48974 13970 49026
rect 14478 48974 14530 49026
rect 15710 48974 15762 49026
rect 16270 48974 16322 49026
rect 16942 48974 16994 49026
rect 17502 48974 17554 49026
rect 19182 48974 19234 49026
rect 19966 48974 20018 49026
rect 21758 48974 21810 49026
rect 22318 48974 22370 49026
rect 23550 48974 23602 49026
rect 24110 48974 24162 49026
rect 26238 48974 26290 49026
rect 27246 48974 27298 49026
rect 28030 48974 28082 49026
rect 28366 48974 28418 49026
rect 28702 48974 28754 49026
rect 29150 48974 29202 49026
rect 29374 48974 29426 49026
rect 33406 48974 33458 49026
rect 37550 48974 37602 49026
rect 38446 48974 38498 49026
rect 39454 48974 39506 49026
rect 39566 48974 39618 49026
rect 40798 48974 40850 49026
rect 41022 48974 41074 49026
rect 43822 48974 43874 49026
rect 46174 48974 46226 49026
rect 47182 48974 47234 49026
rect 53006 48974 53058 49026
rect 53230 48974 53282 49026
rect 54238 48974 54290 49026
rect 54686 48974 54738 49026
rect 55582 48974 55634 49026
rect 8206 48862 8258 48914
rect 10894 48862 10946 48914
rect 14030 48862 14082 48914
rect 17726 48862 17778 48914
rect 22990 48862 23042 48914
rect 27358 48862 27410 48914
rect 29822 48862 29874 48914
rect 31950 48862 32002 48914
rect 37886 48862 37938 48914
rect 38334 48862 38386 48914
rect 38558 48862 38610 48914
rect 39902 48862 39954 48914
rect 43598 48862 43650 48914
rect 44158 48862 44210 48914
rect 45614 48862 45666 48914
rect 45838 48862 45890 48914
rect 46398 48862 46450 48914
rect 46734 48862 46786 48914
rect 51662 48862 51714 48914
rect 51774 48862 51826 48914
rect 4734 48750 4786 48802
rect 11118 48750 11170 48802
rect 15262 48750 15314 48802
rect 27582 48750 27634 48802
rect 27694 48750 27746 48802
rect 27918 48750 27970 48802
rect 28478 48750 28530 48802
rect 29598 48750 29650 48802
rect 30270 48750 30322 48802
rect 31278 48750 31330 48802
rect 31502 48750 31554 48802
rect 31614 48750 31666 48802
rect 31726 48750 31778 48802
rect 32398 48750 32450 48802
rect 32622 48750 32674 48802
rect 32846 48750 32898 48802
rect 34750 48750 34802 48802
rect 40462 48750 40514 48802
rect 44942 48750 44994 48802
rect 45502 48750 45554 48802
rect 47742 48750 47794 48802
rect 51998 48750 52050 48802
rect 52782 48750 52834 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 8094 48414 8146 48466
rect 11566 48414 11618 48466
rect 23326 48414 23378 48466
rect 24222 48414 24274 48466
rect 26798 48414 26850 48466
rect 27470 48414 27522 48466
rect 29374 48414 29426 48466
rect 29822 48414 29874 48466
rect 33070 48414 33122 48466
rect 34526 48414 34578 48466
rect 37102 48414 37154 48466
rect 8990 48302 9042 48354
rect 24670 48302 24722 48354
rect 26126 48302 26178 48354
rect 27582 48302 27634 48354
rect 27694 48302 27746 48354
rect 30606 48302 30658 48354
rect 31502 48302 31554 48354
rect 4286 48190 4338 48242
rect 7982 48190 8034 48242
rect 8766 48190 8818 48242
rect 9886 48190 9938 48242
rect 10446 48190 10498 48242
rect 11230 48190 11282 48242
rect 11342 48190 11394 48242
rect 12462 48190 12514 48242
rect 13470 48190 13522 48242
rect 14814 48190 14866 48242
rect 15262 48190 15314 48242
rect 15598 48190 15650 48242
rect 18622 48190 18674 48242
rect 19294 48190 19346 48242
rect 20078 48190 20130 48242
rect 21086 48190 21138 48242
rect 22318 48190 22370 48242
rect 22878 48190 22930 48242
rect 25790 48190 25842 48242
rect 26798 48190 26850 48242
rect 27246 48190 27298 48242
rect 39006 48414 39058 48466
rect 40126 48414 40178 48466
rect 41022 48414 41074 48466
rect 43486 48414 43538 48466
rect 44270 48414 44322 48466
rect 44830 48414 44882 48466
rect 46174 48414 46226 48466
rect 47070 48414 47122 48466
rect 33630 48302 33682 48354
rect 35086 48302 35138 48354
rect 37774 48302 37826 48354
rect 37998 48302 38050 48354
rect 40910 48302 40962 48354
rect 45166 48302 45218 48354
rect 49422 48302 49474 48354
rect 50878 48302 50930 48354
rect 53230 48302 53282 48354
rect 30270 48190 30322 48242
rect 33070 48190 33122 48242
rect 33518 48190 33570 48242
rect 34414 48190 34466 48242
rect 34974 48190 35026 48242
rect 35982 48190 36034 48242
rect 38222 48190 38274 48242
rect 39902 48190 39954 48242
rect 41246 48190 41298 48242
rect 43822 48190 43874 48242
rect 45502 48190 45554 48242
rect 46062 48190 46114 48242
rect 47406 48190 47458 48242
rect 48974 48190 49026 48242
rect 49198 48190 49250 48242
rect 50318 48190 50370 48242
rect 52110 48190 52162 48242
rect 52446 48190 52498 48242
rect 52670 48190 52722 48242
rect 7646 48078 7698 48130
rect 11566 48078 11618 48130
rect 18510 48078 18562 48130
rect 25454 48078 25506 48130
rect 28030 48078 28082 48130
rect 28366 48078 28418 48130
rect 28590 48078 28642 48130
rect 31054 48078 31106 48130
rect 32062 48078 32114 48130
rect 32622 48078 32674 48130
rect 33182 48078 33234 48130
rect 35534 48078 35586 48130
rect 35758 48078 35810 48130
rect 37662 48078 37714 48130
rect 39454 48078 39506 48130
rect 41694 48078 41746 48130
rect 44158 48078 44210 48130
rect 46734 48078 46786 48130
rect 47742 48078 47794 48130
rect 50094 48078 50146 48130
rect 52558 48078 52610 48130
rect 53118 48078 53170 48130
rect 1934 47966 1986 48018
rect 13470 47966 13522 48018
rect 20638 47966 20690 48018
rect 28926 47966 28978 48018
rect 38670 47966 38722 48018
rect 40238 47966 40290 48018
rect 47854 47966 47906 48018
rect 49534 47966 49586 48018
rect 53006 47966 53058 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 7422 47630 7474 47682
rect 19182 47630 19234 47682
rect 30494 47630 30546 47682
rect 31726 47630 31778 47682
rect 35758 47630 35810 47682
rect 47406 47630 47458 47682
rect 47854 47630 47906 47682
rect 9550 47518 9602 47570
rect 10670 47518 10722 47570
rect 11454 47518 11506 47570
rect 14926 47518 14978 47570
rect 17054 47518 17106 47570
rect 19854 47518 19906 47570
rect 20750 47518 20802 47570
rect 22430 47518 22482 47570
rect 24670 47518 24722 47570
rect 25566 47518 25618 47570
rect 27246 47518 27298 47570
rect 27694 47518 27746 47570
rect 28478 47518 28530 47570
rect 29598 47518 29650 47570
rect 31390 47518 31442 47570
rect 32846 47518 32898 47570
rect 39342 47518 39394 47570
rect 41246 47518 41298 47570
rect 46734 47518 46786 47570
rect 52894 47518 52946 47570
rect 53678 47518 53730 47570
rect 11006 47406 11058 47458
rect 12350 47406 12402 47458
rect 12910 47406 12962 47458
rect 13470 47406 13522 47458
rect 15822 47406 15874 47458
rect 16382 47406 16434 47458
rect 17278 47406 17330 47458
rect 18062 47406 18114 47458
rect 18286 47406 18338 47458
rect 19294 47406 19346 47458
rect 20190 47406 20242 47458
rect 21310 47406 21362 47458
rect 22766 47406 22818 47458
rect 23774 47406 23826 47458
rect 25118 47406 25170 47458
rect 25342 47406 25394 47458
rect 26014 47406 26066 47458
rect 28254 47406 28306 47458
rect 31166 47406 31218 47458
rect 31950 47406 32002 47458
rect 33406 47406 33458 47458
rect 33630 47406 33682 47458
rect 35310 47406 35362 47458
rect 37214 47406 37266 47458
rect 37438 47406 37490 47458
rect 37662 47406 37714 47458
rect 38110 47406 38162 47458
rect 40238 47406 40290 47458
rect 40798 47406 40850 47458
rect 41918 47406 41970 47458
rect 43710 47406 43762 47458
rect 45166 47406 45218 47458
rect 45390 47406 45442 47458
rect 45502 47406 45554 47458
rect 45950 47406 46002 47458
rect 46958 47406 47010 47458
rect 47182 47406 47234 47458
rect 49758 47406 49810 47458
rect 50206 47406 50258 47458
rect 53118 47406 53170 47458
rect 7310 47294 7362 47346
rect 14030 47294 14082 47346
rect 16718 47294 16770 47346
rect 21422 47294 21474 47346
rect 22318 47294 22370 47346
rect 22654 47294 22706 47346
rect 23214 47294 23266 47346
rect 25678 47294 25730 47346
rect 26350 47294 26402 47346
rect 26574 47294 26626 47346
rect 28030 47294 28082 47346
rect 28590 47294 28642 47346
rect 29150 47294 29202 47346
rect 29374 47294 29426 47346
rect 29710 47294 29762 47346
rect 30382 47294 30434 47346
rect 33742 47294 33794 47346
rect 34190 47294 34242 47346
rect 35086 47294 35138 47346
rect 40910 47294 40962 47346
rect 41694 47294 41746 47346
rect 44270 47294 44322 47346
rect 48078 47294 48130 47346
rect 50766 47294 50818 47346
rect 8654 47182 8706 47234
rect 9214 47182 9266 47234
rect 9998 47182 10050 47234
rect 12014 47182 12066 47234
rect 21870 47182 21922 47234
rect 36094 47182 36146 47234
rect 37886 47182 37938 47234
rect 38222 47182 38274 47234
rect 39230 47182 39282 47234
rect 51774 47182 51826 47234
rect 58158 47182 58210 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 11678 46846 11730 46898
rect 13134 46846 13186 46898
rect 13582 46846 13634 46898
rect 16046 46846 16098 46898
rect 16830 46846 16882 46898
rect 18062 46846 18114 46898
rect 20414 46846 20466 46898
rect 20974 46846 21026 46898
rect 29486 46846 29538 46898
rect 33182 46846 33234 46898
rect 35086 46846 35138 46898
rect 38782 46846 38834 46898
rect 39118 46846 39170 46898
rect 40126 46846 40178 46898
rect 40350 46846 40402 46898
rect 45838 46846 45890 46898
rect 50990 46846 51042 46898
rect 53678 46846 53730 46898
rect 6750 46734 6802 46786
rect 8766 46734 8818 46786
rect 9998 46734 10050 46786
rect 10558 46734 10610 46786
rect 11230 46734 11282 46786
rect 11902 46734 11954 46786
rect 14030 46734 14082 46786
rect 14478 46734 14530 46786
rect 14590 46734 14642 46786
rect 16270 46734 16322 46786
rect 21310 46734 21362 46786
rect 27470 46734 27522 46786
rect 29598 46734 29650 46786
rect 29822 46734 29874 46786
rect 30158 46734 30210 46786
rect 34974 46734 35026 46786
rect 35534 46734 35586 46786
rect 36318 46734 36370 46786
rect 39902 46734 39954 46786
rect 41022 46734 41074 46786
rect 44046 46734 44098 46786
rect 45502 46734 45554 46786
rect 48750 46734 48802 46786
rect 49086 46734 49138 46786
rect 50318 46734 50370 46786
rect 52782 46734 52834 46786
rect 7086 46622 7138 46674
rect 9774 46622 9826 46674
rect 10334 46622 10386 46674
rect 12014 46622 12066 46674
rect 12462 46622 12514 46674
rect 17390 46622 17442 46674
rect 17950 46622 18002 46674
rect 18174 46622 18226 46674
rect 18286 46622 18338 46674
rect 18734 46622 18786 46674
rect 18958 46622 19010 46674
rect 19742 46622 19794 46674
rect 20190 46622 20242 46674
rect 22206 46622 22258 46674
rect 22430 46622 22482 46674
rect 22878 46622 22930 46674
rect 23774 46622 23826 46674
rect 27918 46622 27970 46674
rect 28926 46622 28978 46674
rect 29262 46622 29314 46674
rect 30270 46622 30322 46674
rect 32510 46622 32562 46674
rect 35198 46622 35250 46674
rect 35982 46622 36034 46674
rect 36990 46622 37042 46674
rect 40238 46622 40290 46674
rect 40910 46622 40962 46674
rect 41806 46622 41858 46674
rect 42478 46622 42530 46674
rect 42926 46622 42978 46674
rect 44942 46622 44994 46674
rect 45166 46622 45218 46674
rect 46062 46622 46114 46674
rect 48862 46622 48914 46674
rect 49534 46622 49586 46674
rect 50206 46622 50258 46674
rect 50542 46622 50594 46674
rect 51774 46622 51826 46674
rect 51998 46622 52050 46674
rect 52222 46622 52274 46674
rect 52334 46622 52386 46674
rect 52670 46622 52722 46674
rect 53566 46622 53618 46674
rect 11566 46510 11618 46562
rect 16494 46510 16546 46562
rect 20302 46510 20354 46562
rect 21870 46510 21922 46562
rect 24110 46510 24162 46562
rect 25230 46510 25282 46562
rect 26574 46510 26626 46562
rect 27022 46510 27074 46562
rect 28366 46510 28418 46562
rect 31726 46510 31778 46562
rect 34638 46510 34690 46562
rect 36654 46510 36706 46562
rect 36766 46510 36818 46562
rect 37998 46510 38050 46562
rect 38446 46510 38498 46562
rect 41470 46510 41522 46562
rect 45390 46510 45442 46562
rect 49310 46510 49362 46562
rect 49982 46510 50034 46562
rect 8542 46398 8594 46450
rect 8878 46398 8930 46450
rect 14254 46398 14306 46450
rect 14814 46398 14866 46450
rect 15038 46398 15090 46450
rect 17614 46398 17666 46450
rect 19406 46398 19458 46450
rect 20638 46398 20690 46450
rect 21086 46398 21138 46450
rect 21534 46398 21586 46450
rect 23998 46398 24050 46450
rect 25454 46398 25506 46450
rect 25790 46398 25842 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 15710 46062 15762 46114
rect 17614 46062 17666 46114
rect 32846 46062 32898 46114
rect 33854 46062 33906 46114
rect 34638 46062 34690 46114
rect 41246 46062 41298 46114
rect 10334 45950 10386 46002
rect 16382 45950 16434 46002
rect 17502 45950 17554 46002
rect 18734 45950 18786 46002
rect 20302 45950 20354 46002
rect 23102 45950 23154 46002
rect 23886 45950 23938 46002
rect 24782 45950 24834 46002
rect 26238 45950 26290 46002
rect 27358 45950 27410 46002
rect 28590 45950 28642 46002
rect 30046 45950 30098 46002
rect 33854 45950 33906 46002
rect 47966 45950 48018 46002
rect 6078 45838 6130 45890
rect 7198 45838 7250 45890
rect 7646 45838 7698 45890
rect 8094 45838 8146 45890
rect 8878 45838 8930 45890
rect 9550 45838 9602 45890
rect 10110 45838 10162 45890
rect 11790 45838 11842 45890
rect 14142 45838 14194 45890
rect 14366 45838 14418 45890
rect 15486 45838 15538 45890
rect 15598 45838 15650 45890
rect 15934 45838 15986 45890
rect 18958 45838 19010 45890
rect 19182 45838 19234 45890
rect 21310 45838 21362 45890
rect 21870 45838 21922 45890
rect 23774 45838 23826 45890
rect 24670 45838 24722 45890
rect 25678 45838 25730 45890
rect 26574 45838 26626 45890
rect 27694 45838 27746 45890
rect 30158 45838 30210 45890
rect 30382 45838 30434 45890
rect 31278 45838 31330 45890
rect 31502 45838 31554 45890
rect 32286 45838 32338 45890
rect 32398 45838 32450 45890
rect 32734 45838 32786 45890
rect 35422 45838 35474 45890
rect 38558 45838 38610 45890
rect 41582 45838 41634 45890
rect 44942 45838 44994 45890
rect 45278 45838 45330 45890
rect 46062 45838 46114 45890
rect 47406 45838 47458 45890
rect 6302 45726 6354 45778
rect 8766 45726 8818 45778
rect 10446 45726 10498 45778
rect 13470 45726 13522 45778
rect 17838 45726 17890 45778
rect 19742 45726 19794 45778
rect 20190 45726 20242 45778
rect 20526 45726 20578 45778
rect 20750 45726 20802 45778
rect 21982 45726 22034 45778
rect 24110 45726 24162 45778
rect 24446 45726 24498 45778
rect 27022 45726 27074 45778
rect 27358 45726 27410 45778
rect 29150 45726 29202 45778
rect 29262 45726 29314 45778
rect 30494 45726 30546 45778
rect 34862 45726 34914 45778
rect 39006 45726 39058 45778
rect 39230 45726 39282 45778
rect 45502 45726 45554 45778
rect 48750 45726 48802 45778
rect 49646 45726 49698 45778
rect 6638 45614 6690 45666
rect 9438 45614 9490 45666
rect 12910 45614 12962 45666
rect 21534 45614 21586 45666
rect 23438 45614 23490 45666
rect 25118 45614 25170 45666
rect 29486 45614 29538 45666
rect 34302 45614 34354 45666
rect 38782 45614 38834 45666
rect 41358 45614 41410 45666
rect 48414 45614 48466 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 13246 45278 13298 45330
rect 17502 45278 17554 45330
rect 17614 45278 17666 45330
rect 18734 45278 18786 45330
rect 21758 45278 21810 45330
rect 22990 45278 23042 45330
rect 23438 45278 23490 45330
rect 23886 45278 23938 45330
rect 24670 45278 24722 45330
rect 25342 45278 25394 45330
rect 25790 45278 25842 45330
rect 28926 45278 28978 45330
rect 31278 45278 31330 45330
rect 34414 45278 34466 45330
rect 53790 45278 53842 45330
rect 10446 45166 10498 45218
rect 11678 45166 11730 45218
rect 14030 45166 14082 45218
rect 19966 45166 20018 45218
rect 20190 45166 20242 45218
rect 20750 45166 20802 45218
rect 24446 45166 24498 45218
rect 24782 45166 24834 45218
rect 27806 45166 27858 45218
rect 29486 45166 29538 45218
rect 29710 45166 29762 45218
rect 30606 45166 30658 45218
rect 31390 45166 31442 45218
rect 33070 45166 33122 45218
rect 33406 45166 33458 45218
rect 34078 45166 34130 45218
rect 34638 45166 34690 45218
rect 40014 45166 40066 45218
rect 42030 45166 42082 45218
rect 45054 45166 45106 45218
rect 45166 45166 45218 45218
rect 45726 45166 45778 45218
rect 47742 45166 47794 45218
rect 48974 45166 49026 45218
rect 49310 45166 49362 45218
rect 53566 45166 53618 45218
rect 55918 45166 55970 45218
rect 7310 45054 7362 45106
rect 10110 45054 10162 45106
rect 11790 45054 11842 45106
rect 12910 45054 12962 45106
rect 13022 45054 13074 45106
rect 13358 45054 13410 45106
rect 19854 45054 19906 45106
rect 20526 45054 20578 45106
rect 24110 45054 24162 45106
rect 26686 45054 26738 45106
rect 27022 45054 27074 45106
rect 27918 45054 27970 45106
rect 28478 45054 28530 45106
rect 28702 45054 28754 45106
rect 28814 45054 28866 45106
rect 29150 45054 29202 45106
rect 30718 45054 30770 45106
rect 31166 45054 31218 45106
rect 32510 45054 32562 45106
rect 34302 45054 34354 45106
rect 35310 45054 35362 45106
rect 35534 45054 35586 45106
rect 36206 45054 36258 45106
rect 40350 45054 40402 45106
rect 41358 45054 41410 45106
rect 42142 45054 42194 45106
rect 45278 45054 45330 45106
rect 46846 45054 46898 45106
rect 47070 45054 47122 45106
rect 48750 45054 48802 45106
rect 50318 45054 50370 45106
rect 50990 45054 51042 45106
rect 54574 45054 54626 45106
rect 55246 45054 55298 45106
rect 55582 45054 55634 45106
rect 7870 44942 7922 44994
rect 14142 44942 14194 44994
rect 14926 44942 14978 44994
rect 15262 44942 15314 44994
rect 15710 44942 15762 44994
rect 16382 44942 16434 44994
rect 16830 44942 16882 44994
rect 18286 44942 18338 44994
rect 19070 44942 19122 44994
rect 19518 44942 19570 44994
rect 21198 44942 21250 44994
rect 22094 44942 22146 44994
rect 26238 44942 26290 44994
rect 28030 44942 28082 44994
rect 29598 44942 29650 44994
rect 38334 44942 38386 44994
rect 41806 44942 41858 44994
rect 46622 44942 46674 44994
rect 49982 44942 50034 44994
rect 50766 44942 50818 44994
rect 53902 44942 53954 44994
rect 54350 44942 54402 44994
rect 13806 44830 13858 44882
rect 17726 44830 17778 44882
rect 36430 44830 36482 44882
rect 40350 44830 40402 44882
rect 47294 44830 47346 44882
rect 51214 44830 51266 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 7534 44494 7586 44546
rect 14814 44494 14866 44546
rect 19294 44494 19346 44546
rect 24894 44494 24946 44546
rect 29262 44494 29314 44546
rect 30046 44494 30098 44546
rect 43374 44494 43426 44546
rect 43486 44494 43538 44546
rect 46734 44494 46786 44546
rect 46958 44494 47010 44546
rect 47406 44494 47458 44546
rect 47518 44494 47570 44546
rect 16718 44382 16770 44434
rect 16942 44382 16994 44434
rect 18846 44382 18898 44434
rect 22318 44382 22370 44434
rect 23998 44382 24050 44434
rect 28590 44382 28642 44434
rect 32622 44382 32674 44434
rect 34526 44382 34578 44434
rect 37886 44382 37938 44434
rect 38222 44382 38274 44434
rect 39230 44382 39282 44434
rect 39342 44382 39394 44434
rect 41358 44382 41410 44434
rect 49310 44382 49362 44434
rect 50878 44382 50930 44434
rect 51326 44382 51378 44434
rect 53678 44382 53730 44434
rect 54686 44382 54738 44434
rect 57934 44382 57986 44434
rect 9998 44270 10050 44322
rect 12910 44270 12962 44322
rect 15710 44270 15762 44322
rect 16606 44270 16658 44322
rect 17278 44270 17330 44322
rect 18510 44270 18562 44322
rect 19070 44270 19122 44322
rect 19854 44270 19906 44322
rect 21310 44270 21362 44322
rect 21870 44270 21922 44322
rect 23886 44270 23938 44322
rect 24110 44270 24162 44322
rect 24558 44270 24610 44322
rect 25006 44270 25058 44322
rect 26462 44270 26514 44322
rect 26798 44270 26850 44322
rect 29486 44270 29538 44322
rect 29710 44270 29762 44322
rect 30606 44270 30658 44322
rect 31838 44270 31890 44322
rect 32286 44270 32338 44322
rect 32846 44270 32898 44322
rect 33966 44270 34018 44322
rect 34974 44270 35026 44322
rect 35982 44270 36034 44322
rect 37550 44270 37602 44322
rect 39006 44270 39058 44322
rect 39678 44270 39730 44322
rect 40798 44270 40850 44322
rect 41022 44270 41074 44322
rect 41246 44270 41298 44322
rect 41470 44270 41522 44322
rect 42702 44270 42754 44322
rect 43150 44270 43202 44322
rect 45054 44270 45106 44322
rect 45390 44270 45442 44322
rect 45838 44270 45890 44322
rect 47294 44270 47346 44322
rect 48862 44270 48914 44322
rect 50654 44270 50706 44322
rect 53790 44270 53842 44322
rect 54574 44270 54626 44322
rect 55918 44270 55970 44322
rect 7310 44158 7362 44210
rect 14478 44158 14530 44210
rect 17614 44158 17666 44210
rect 19966 44158 20018 44210
rect 20526 44158 20578 44210
rect 25342 44158 25394 44210
rect 29822 44158 29874 44210
rect 31054 44158 31106 44210
rect 31278 44158 31330 44210
rect 33070 44158 33122 44210
rect 33854 44158 33906 44210
rect 34526 44158 34578 44210
rect 35646 44158 35698 44210
rect 38782 44158 38834 44210
rect 54910 44158 54962 44210
rect 7870 44046 7922 44098
rect 10110 44046 10162 44098
rect 10334 44046 10386 44098
rect 12350 44046 12402 44098
rect 13582 44046 13634 44098
rect 14030 44046 14082 44098
rect 14702 44046 14754 44098
rect 15150 44046 15202 44098
rect 20190 44046 20242 44098
rect 23102 44046 23154 44098
rect 23550 44046 23602 44098
rect 30942 44046 30994 44098
rect 35758 44046 35810 44098
rect 36318 44046 36370 44098
rect 43486 44046 43538 44098
rect 44830 44046 44882 44098
rect 44942 44046 44994 44098
rect 46062 44046 46114 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 6974 43710 7026 43762
rect 8094 43710 8146 43762
rect 29934 43710 29986 43762
rect 33406 43710 33458 43762
rect 33742 43710 33794 43762
rect 34414 43710 34466 43762
rect 41246 43710 41298 43762
rect 46734 43710 46786 43762
rect 49870 43710 49922 43762
rect 54126 43710 54178 43762
rect 7646 43598 7698 43650
rect 14366 43598 14418 43650
rect 14926 43598 14978 43650
rect 18398 43598 18450 43650
rect 21086 43598 21138 43650
rect 23214 43598 23266 43650
rect 23438 43598 23490 43650
rect 24334 43598 24386 43650
rect 27022 43598 27074 43650
rect 29038 43598 29090 43650
rect 29150 43598 29202 43650
rect 30830 43598 30882 43650
rect 31390 43598 31442 43650
rect 34638 43598 34690 43650
rect 36654 43598 36706 43650
rect 36766 43598 36818 43650
rect 51438 43598 51490 43650
rect 53118 43598 53170 43650
rect 53902 43598 53954 43650
rect 56590 43598 56642 43650
rect 6638 43486 6690 43538
rect 7422 43486 7474 43538
rect 7534 43486 7586 43538
rect 9550 43486 9602 43538
rect 11118 43486 11170 43538
rect 12350 43486 12402 43538
rect 13358 43486 13410 43538
rect 13918 43486 13970 43538
rect 14814 43486 14866 43538
rect 16158 43486 16210 43538
rect 17726 43486 17778 43538
rect 18174 43486 18226 43538
rect 18958 43486 19010 43538
rect 19518 43486 19570 43538
rect 20414 43486 20466 43538
rect 20974 43486 21026 43538
rect 21870 43486 21922 43538
rect 23774 43486 23826 43538
rect 25342 43486 25394 43538
rect 25566 43486 25618 43538
rect 26574 43486 26626 43538
rect 28030 43486 28082 43538
rect 29598 43486 29650 43538
rect 30382 43486 30434 43538
rect 34862 43486 34914 43538
rect 36430 43486 36482 43538
rect 37774 43486 37826 43538
rect 40910 43486 40962 43538
rect 42590 43486 42642 43538
rect 43710 43486 43762 43538
rect 44382 43486 44434 43538
rect 45278 43486 45330 43538
rect 49086 43486 49138 43538
rect 51326 43486 51378 43538
rect 51662 43486 51714 43538
rect 52222 43486 52274 43538
rect 53454 43486 53506 43538
rect 54798 43486 54850 43538
rect 55470 43486 55522 43538
rect 56814 43486 56866 43538
rect 10334 43374 10386 43426
rect 15710 43374 15762 43426
rect 16494 43374 16546 43426
rect 17390 43374 17442 43426
rect 21646 43374 21698 43426
rect 22766 43374 22818 43426
rect 27694 43374 27746 43426
rect 34750 43374 34802 43426
rect 38446 43374 38498 43426
rect 38558 43374 38610 43426
rect 46174 43374 46226 43426
rect 49310 43374 49362 43426
rect 52334 43374 52386 43426
rect 54014 43374 54066 43426
rect 54574 43374 54626 43426
rect 11118 43262 11170 43314
rect 11454 43262 11506 43314
rect 14926 43262 14978 43314
rect 23102 43262 23154 43314
rect 26462 43262 26514 43314
rect 28254 43262 28306 43314
rect 28590 43262 28642 43314
rect 29038 43262 29090 43314
rect 37214 43262 37266 43314
rect 45278 43262 45330 43314
rect 49422 43262 49474 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 16606 42926 16658 42978
rect 18734 42926 18786 42978
rect 28030 42926 28082 42978
rect 29598 42926 29650 42978
rect 30718 42926 30770 42978
rect 36318 42926 36370 42978
rect 45838 42926 45890 42978
rect 57934 42926 57986 42978
rect 1710 42814 1762 42866
rect 7646 42814 7698 42866
rect 12126 42814 12178 42866
rect 12686 42814 12738 42866
rect 18286 42814 18338 42866
rect 19518 42814 19570 42866
rect 21534 42814 21586 42866
rect 26574 42814 26626 42866
rect 27470 42814 27522 42866
rect 29822 42814 29874 42866
rect 34414 42814 34466 42866
rect 37774 42814 37826 42866
rect 38446 42814 38498 42866
rect 42926 42814 42978 42866
rect 45390 42814 45442 42866
rect 51214 42814 51266 42866
rect 52782 42814 52834 42866
rect 53678 42814 53730 42866
rect 7310 42702 7362 42754
rect 7870 42702 7922 42754
rect 10334 42702 10386 42754
rect 13806 42702 13858 42754
rect 15038 42702 15090 42754
rect 16046 42702 16098 42754
rect 17614 42702 17666 42754
rect 18734 42702 18786 42754
rect 19742 42702 19794 42754
rect 20526 42702 20578 42754
rect 21310 42702 21362 42754
rect 22318 42702 22370 42754
rect 22990 42702 23042 42754
rect 24446 42702 24498 42754
rect 25902 42702 25954 42754
rect 26798 42702 26850 42754
rect 27582 42702 27634 42754
rect 28702 42702 28754 42754
rect 29038 42702 29090 42754
rect 30382 42702 30434 42754
rect 31838 42702 31890 42754
rect 32398 42702 32450 42754
rect 34302 42702 34354 42754
rect 36094 42702 36146 42754
rect 37438 42702 37490 42754
rect 37550 42702 37602 42754
rect 38558 42702 38610 42754
rect 41358 42702 41410 42754
rect 41918 42702 41970 42754
rect 42254 42702 42306 42754
rect 44942 42702 44994 42754
rect 45502 42702 45554 42754
rect 47966 42702 48018 42754
rect 48190 42702 48242 42754
rect 48414 42702 48466 42754
rect 49422 42702 49474 42754
rect 53006 42702 53058 42754
rect 56030 42702 56082 42754
rect 8318 42590 8370 42642
rect 9774 42590 9826 42642
rect 10894 42590 10946 42642
rect 16270 42590 16322 42642
rect 19406 42590 19458 42642
rect 24894 42590 24946 42642
rect 26014 42590 26066 42642
rect 29374 42590 29426 42642
rect 30046 42590 30098 42642
rect 31502 42590 31554 42642
rect 32510 42590 32562 42642
rect 32734 42590 32786 42642
rect 35534 42590 35586 42642
rect 37886 42590 37938 42642
rect 38222 42590 38274 42642
rect 42590 42590 42642 42642
rect 49982 42590 50034 42642
rect 9214 42478 9266 42530
rect 21870 42478 21922 42530
rect 24110 42478 24162 42530
rect 30158 42478 30210 42530
rect 30606 42478 30658 42530
rect 31166 42478 31218 42530
rect 31614 42478 31666 42530
rect 39006 42478 39058 42530
rect 48862 42478 48914 42530
rect 50878 42478 50930 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 8542 42142 8594 42194
rect 13918 42142 13970 42194
rect 21646 42142 21698 42194
rect 27918 42142 27970 42194
rect 30270 42142 30322 42194
rect 30830 42142 30882 42194
rect 33182 42142 33234 42194
rect 33742 42142 33794 42194
rect 41358 42142 41410 42194
rect 42366 42142 42418 42194
rect 46510 42142 46562 42194
rect 49086 42142 49138 42194
rect 51550 42142 51602 42194
rect 51774 42142 51826 42194
rect 52558 42142 52610 42194
rect 10782 42030 10834 42082
rect 12574 42030 12626 42082
rect 13470 42030 13522 42082
rect 15486 42030 15538 42082
rect 19630 42030 19682 42082
rect 19966 42030 20018 42082
rect 20750 42030 20802 42082
rect 22990 42030 23042 42082
rect 23662 42030 23714 42082
rect 25566 42030 25618 42082
rect 27470 42030 27522 42082
rect 28142 42030 28194 42082
rect 28926 42030 28978 42082
rect 29150 42030 29202 42082
rect 31054 42030 31106 42082
rect 34862 42030 34914 42082
rect 35086 42030 35138 42082
rect 35646 42030 35698 42082
rect 47518 42030 47570 42082
rect 49310 42030 49362 42082
rect 11342 41918 11394 41970
rect 12126 41918 12178 41970
rect 12462 41918 12514 41970
rect 14590 41918 14642 41970
rect 14926 41918 14978 41970
rect 17390 41918 17442 41970
rect 18286 41918 18338 41970
rect 19406 41918 19458 41970
rect 19742 41918 19794 41970
rect 21422 41918 21474 41970
rect 21534 41918 21586 41970
rect 21870 41918 21922 41970
rect 22654 41918 22706 41970
rect 22878 41918 22930 41970
rect 23886 41918 23938 41970
rect 25342 41918 25394 41970
rect 26462 41918 26514 41970
rect 27358 41918 27410 41970
rect 28478 41918 28530 41970
rect 29374 41918 29426 41970
rect 29822 41918 29874 41970
rect 30494 41918 30546 41970
rect 31166 41918 31218 41970
rect 34190 41918 34242 41970
rect 34638 41918 34690 41970
rect 35198 41918 35250 41970
rect 35870 41918 35922 41970
rect 39790 41918 39842 41970
rect 42142 41918 42194 41970
rect 42478 41918 42530 41970
rect 45278 41918 45330 41970
rect 45726 41918 45778 41970
rect 45950 41918 46002 41970
rect 46286 41918 46338 41970
rect 47294 41918 47346 41970
rect 47742 41918 47794 41970
rect 47854 41918 47906 41970
rect 48750 41918 48802 41970
rect 49198 41918 49250 41970
rect 49758 41918 49810 41970
rect 50094 41918 50146 41970
rect 51214 41918 51266 41970
rect 51886 41918 51938 41970
rect 52446 41918 52498 41970
rect 52782 41918 52834 41970
rect 7982 41806 8034 41858
rect 17950 41806 18002 41858
rect 22094 41806 22146 41858
rect 25678 41806 25730 41858
rect 29262 41806 29314 41858
rect 34974 41806 35026 41858
rect 40238 41806 40290 41858
rect 41918 41806 41970 41858
rect 44382 41806 44434 41858
rect 44830 41806 44882 41858
rect 50654 41806 50706 41858
rect 8206 41694 8258 41746
rect 18398 41694 18450 41746
rect 22318 41694 22370 41746
rect 29598 41694 29650 41746
rect 30270 41694 30322 41746
rect 33630 41694 33682 41746
rect 34302 41694 34354 41746
rect 46174 41694 46226 41746
rect 47070 41694 47122 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 17166 41358 17218 41410
rect 21422 41358 21474 41410
rect 26014 41358 26066 41410
rect 37550 41358 37602 41410
rect 42030 41358 42082 41410
rect 47294 41358 47346 41410
rect 1710 41246 1762 41298
rect 8542 41246 8594 41298
rect 11678 41246 11730 41298
rect 18846 41246 18898 41298
rect 20862 41246 20914 41298
rect 22542 41246 22594 41298
rect 22766 41246 22818 41298
rect 23438 41246 23490 41298
rect 24222 41246 24274 41298
rect 27806 41246 27858 41298
rect 30046 41246 30098 41298
rect 34078 41246 34130 41298
rect 34638 41246 34690 41298
rect 40462 41246 40514 41298
rect 42590 41246 42642 41298
rect 46622 41246 46674 41298
rect 48078 41246 48130 41298
rect 49086 41246 49138 41298
rect 52894 41246 52946 41298
rect 57934 41246 57986 41298
rect 7086 41134 7138 41186
rect 8318 41134 8370 41186
rect 8990 41134 9042 41186
rect 10558 41134 10610 41186
rect 11454 41134 11506 41186
rect 12686 41134 12738 41186
rect 13470 41134 13522 41186
rect 14366 41134 14418 41186
rect 14814 41134 14866 41186
rect 16046 41134 16098 41186
rect 17166 41134 17218 41186
rect 17390 41134 17442 41186
rect 17950 41134 18002 41186
rect 18174 41134 18226 41186
rect 18958 41134 19010 41186
rect 21534 41134 21586 41186
rect 22318 41134 22370 41186
rect 22878 41134 22930 41186
rect 24558 41134 24610 41186
rect 25454 41134 25506 41186
rect 27022 41134 27074 41186
rect 29598 41134 29650 41186
rect 30606 41134 30658 41186
rect 31502 41134 31554 41186
rect 32622 41134 32674 41186
rect 33630 41134 33682 41186
rect 34414 41134 34466 41186
rect 34750 41134 34802 41186
rect 35086 41134 35138 41186
rect 37214 41134 37266 41186
rect 38782 41134 38834 41186
rect 39230 41134 39282 41186
rect 39678 41134 39730 41186
rect 40910 41134 40962 41186
rect 41694 41134 41746 41186
rect 42926 41134 42978 41186
rect 45614 41134 45666 41186
rect 46398 41134 46450 41186
rect 47518 41134 47570 41186
rect 47854 41134 47906 41186
rect 48638 41134 48690 41186
rect 52670 41134 52722 41186
rect 54574 41134 54626 41186
rect 56030 41134 56082 41186
rect 7310 41022 7362 41074
rect 9214 41022 9266 41074
rect 9662 41022 9714 41074
rect 14254 41022 14306 41074
rect 19630 41022 19682 41074
rect 21422 41022 21474 41074
rect 26238 41022 26290 41074
rect 26686 41022 26738 41074
rect 28702 41022 28754 41074
rect 30830 41022 30882 41074
rect 31166 41022 31218 41074
rect 36990 41022 37042 41074
rect 41134 41022 41186 41074
rect 43486 41022 43538 41074
rect 46734 41022 46786 41074
rect 51326 41022 51378 41074
rect 51550 41022 51602 41074
rect 51774 41022 51826 41074
rect 51886 41022 51938 41074
rect 53006 41022 53058 41074
rect 53342 41022 53394 41074
rect 54350 41022 54402 41074
rect 54462 41022 54514 41074
rect 20078 40910 20130 40962
rect 24782 40910 24834 40962
rect 25678 40910 25730 40962
rect 26126 40910 26178 40962
rect 26798 40910 26850 40962
rect 27358 40910 27410 40962
rect 31502 40910 31554 40962
rect 36542 40910 36594 40962
rect 48190 40910 48242 40962
rect 53454 40910 53506 40962
rect 55022 40910 55074 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 7198 40574 7250 40626
rect 8878 40574 8930 40626
rect 9886 40574 9938 40626
rect 12798 40574 12850 40626
rect 16270 40574 16322 40626
rect 16382 40574 16434 40626
rect 16494 40574 16546 40626
rect 20750 40574 20802 40626
rect 22206 40574 22258 40626
rect 22430 40574 22482 40626
rect 22990 40574 23042 40626
rect 26574 40574 26626 40626
rect 28702 40574 28754 40626
rect 29710 40574 29762 40626
rect 30270 40574 30322 40626
rect 30606 40574 30658 40626
rect 30830 40574 30882 40626
rect 32062 40574 32114 40626
rect 34190 40574 34242 40626
rect 34862 40574 34914 40626
rect 41694 40574 41746 40626
rect 41806 40574 41858 40626
rect 41918 40574 41970 40626
rect 42142 40574 42194 40626
rect 49982 40574 50034 40626
rect 50990 40574 51042 40626
rect 52110 40574 52162 40626
rect 53454 40574 53506 40626
rect 53678 40574 53730 40626
rect 55246 40574 55298 40626
rect 7534 40462 7586 40514
rect 10222 40462 10274 40514
rect 21198 40462 21250 40514
rect 27134 40462 27186 40514
rect 27358 40462 27410 40514
rect 27694 40462 27746 40514
rect 28366 40462 28418 40514
rect 28590 40462 28642 40514
rect 31278 40462 31330 40514
rect 31838 40462 31890 40514
rect 34974 40462 35026 40514
rect 45838 40462 45890 40514
rect 49422 40462 49474 40514
rect 50542 40462 50594 40514
rect 51662 40462 51714 40514
rect 53342 40462 53394 40514
rect 54462 40462 54514 40514
rect 56590 40462 56642 40514
rect 10110 40350 10162 40402
rect 11342 40350 11394 40402
rect 12014 40350 12066 40402
rect 12686 40350 12738 40402
rect 13694 40350 13746 40402
rect 14814 40350 14866 40402
rect 15822 40350 15874 40402
rect 16942 40350 16994 40402
rect 17838 40350 17890 40402
rect 19294 40350 19346 40402
rect 21646 40350 21698 40402
rect 22094 40350 22146 40402
rect 23774 40350 23826 40402
rect 24334 40350 24386 40402
rect 25342 40350 25394 40402
rect 25678 40350 25730 40402
rect 25790 40350 25842 40402
rect 28030 40350 28082 40402
rect 30494 40350 30546 40402
rect 31166 40350 31218 40402
rect 31502 40350 31554 40402
rect 31726 40350 31778 40402
rect 32174 40350 32226 40402
rect 35086 40350 35138 40402
rect 35198 40350 35250 40402
rect 35422 40350 35474 40402
rect 38334 40350 38386 40402
rect 45278 40350 45330 40402
rect 46286 40350 46338 40402
rect 46734 40350 46786 40402
rect 48862 40350 48914 40402
rect 49310 40350 49362 40402
rect 49534 40350 49586 40402
rect 50766 40350 50818 40402
rect 51326 40350 51378 40402
rect 51550 40350 51602 40402
rect 54574 40350 54626 40402
rect 55134 40350 55186 40402
rect 56926 40350 56978 40402
rect 8206 40238 8258 40290
rect 17390 40238 17442 40290
rect 19742 40238 19794 40290
rect 37998 40238 38050 40290
rect 44494 40238 44546 40290
rect 44942 40238 44994 40290
rect 56814 40238 56866 40290
rect 8094 40126 8146 40178
rect 8430 40126 8482 40178
rect 14926 40126 14978 40178
rect 38670 40126 38722 40178
rect 51102 40126 51154 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 9774 39790 9826 39842
rect 11342 39790 11394 39842
rect 22654 39790 22706 39842
rect 23214 39790 23266 39842
rect 23438 39790 23490 39842
rect 29374 39790 29426 39842
rect 29598 39790 29650 39842
rect 37326 39790 37378 39842
rect 37550 39790 37602 39842
rect 37998 39790 38050 39842
rect 38334 39790 38386 39842
rect 42366 39790 42418 39842
rect 49086 39790 49138 39842
rect 49758 39790 49810 39842
rect 54126 39790 54178 39842
rect 12798 39678 12850 39730
rect 19182 39678 19234 39730
rect 20750 39678 20802 39730
rect 22430 39678 22482 39730
rect 23102 39678 23154 39730
rect 24222 39678 24274 39730
rect 25006 39678 25058 39730
rect 26014 39678 26066 39730
rect 28030 39678 28082 39730
rect 31726 39678 31778 39730
rect 33518 39678 33570 39730
rect 35870 39678 35922 39730
rect 49198 39678 49250 39730
rect 49870 39678 49922 39730
rect 57934 39678 57986 39730
rect 6638 39566 6690 39618
rect 7310 39566 7362 39618
rect 7982 39566 8034 39618
rect 8654 39566 8706 39618
rect 9214 39566 9266 39618
rect 9998 39566 10050 39618
rect 10670 39566 10722 39618
rect 11902 39566 11954 39618
rect 13470 39566 13522 39618
rect 14030 39566 14082 39618
rect 14702 39566 14754 39618
rect 15374 39566 15426 39618
rect 16606 39566 16658 39618
rect 16942 39566 16994 39618
rect 19294 39566 19346 39618
rect 21310 39566 21362 39618
rect 21646 39566 21698 39618
rect 21982 39566 22034 39618
rect 22094 39566 22146 39618
rect 22206 39566 22258 39618
rect 23662 39566 23714 39618
rect 24446 39566 24498 39618
rect 27694 39566 27746 39618
rect 27918 39566 27970 39618
rect 29150 39566 29202 39618
rect 32062 39566 32114 39618
rect 34302 39566 34354 39618
rect 34862 39566 34914 39618
rect 35422 39566 35474 39618
rect 37774 39566 37826 39618
rect 39566 39566 39618 39618
rect 42142 39566 42194 39618
rect 45166 39566 45218 39618
rect 45838 39566 45890 39618
rect 46734 39566 46786 39618
rect 48414 39566 48466 39618
rect 48638 39566 48690 39618
rect 51102 39566 51154 39618
rect 56030 39566 56082 39618
rect 6862 39454 6914 39506
rect 8206 39454 8258 39506
rect 14590 39454 14642 39506
rect 19742 39454 19794 39506
rect 25118 39454 25170 39506
rect 29710 39454 29762 39506
rect 32286 39454 32338 39506
rect 35758 39454 35810 39506
rect 45950 39454 46002 39506
rect 48974 39454 49026 39506
rect 49646 39454 49698 39506
rect 50990 39454 51042 39506
rect 54238 39454 54290 39506
rect 1710 39342 1762 39394
rect 7534 39342 7586 39394
rect 15486 39342 15538 39394
rect 24894 39342 24946 39394
rect 28590 39342 28642 39394
rect 35982 39342 36034 39394
rect 39902 39342 39954 39394
rect 42702 39342 42754 39394
rect 44830 39342 44882 39394
rect 46846 39342 46898 39394
rect 54126 39342 54178 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 9550 39006 9602 39058
rect 10782 39006 10834 39058
rect 11678 39006 11730 39058
rect 12574 39006 12626 39058
rect 13470 39006 13522 39058
rect 16270 39006 16322 39058
rect 18398 39006 18450 39058
rect 19182 39006 19234 39058
rect 19518 39006 19570 39058
rect 20750 39006 20802 39058
rect 22206 39006 22258 39058
rect 22430 39006 22482 39058
rect 22654 39006 22706 39058
rect 23998 39006 24050 39058
rect 33406 39006 33458 39058
rect 33854 39006 33906 39058
rect 35198 39006 35250 39058
rect 42590 39006 42642 39058
rect 43598 39006 43650 39058
rect 47854 39006 47906 39058
rect 49646 39006 49698 39058
rect 50094 39006 50146 39058
rect 53230 39006 53282 39058
rect 7646 38894 7698 38946
rect 16830 38894 16882 38946
rect 17838 38894 17890 38946
rect 20862 38894 20914 38946
rect 22878 38894 22930 38946
rect 28478 38894 28530 38946
rect 34862 38894 34914 38946
rect 35758 38894 35810 38946
rect 41806 38894 41858 38946
rect 43038 38894 43090 38946
rect 45614 38894 45666 38946
rect 46286 38894 46338 38946
rect 50542 38894 50594 38946
rect 54798 38894 54850 38946
rect 11342 38782 11394 38834
rect 12238 38782 12290 38834
rect 14030 38782 14082 38834
rect 14814 38782 14866 38834
rect 15262 38782 15314 38834
rect 17950 38782 18002 38834
rect 18286 38782 18338 38834
rect 21870 38782 21922 38834
rect 22990 38782 23042 38834
rect 24110 38782 24162 38834
rect 27806 38782 27858 38834
rect 29262 38782 29314 38834
rect 29486 38782 29538 38834
rect 31726 38782 31778 38834
rect 31950 38782 32002 38834
rect 32286 38782 32338 38834
rect 35534 38782 35586 38834
rect 36094 38782 36146 38834
rect 38558 38782 38610 38834
rect 42142 38782 42194 38834
rect 42478 38782 42530 38834
rect 43262 38782 43314 38834
rect 44718 38782 44770 38834
rect 45054 38782 45106 38834
rect 45166 38782 45218 38834
rect 45950 38782 46002 38834
rect 46398 38782 46450 38834
rect 47294 38782 47346 38834
rect 48974 38782 49026 38834
rect 49198 38782 49250 38834
rect 53118 38782 53170 38834
rect 53454 38782 53506 38834
rect 54126 38782 54178 38834
rect 7870 38670 7922 38722
rect 8430 38670 8482 38722
rect 9998 38670 10050 38722
rect 13134 38670 13186 38722
rect 19966 38670 20018 38722
rect 22318 38670 22370 38722
rect 23998 38670 24050 38722
rect 32510 38670 32562 38722
rect 35982 38670 36034 38722
rect 38334 38670 38386 38722
rect 39230 38670 39282 38722
rect 48750 38670 48802 38722
rect 54014 38670 54066 38722
rect 14590 38558 14642 38610
rect 20638 38558 20690 38610
rect 27694 38558 27746 38610
rect 32398 38558 32450 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 14814 38222 14866 38274
rect 15150 38222 15202 38274
rect 33294 38222 33346 38274
rect 46062 38222 46114 38274
rect 53230 38222 53282 38274
rect 14590 38110 14642 38162
rect 16158 38110 16210 38162
rect 17054 38110 17106 38162
rect 19294 38110 19346 38162
rect 24558 38110 24610 38162
rect 27918 38110 27970 38162
rect 30158 38110 30210 38162
rect 32174 38110 32226 38162
rect 34190 38110 34242 38162
rect 35758 38110 35810 38162
rect 43374 38110 43426 38162
rect 45278 38110 45330 38162
rect 51438 38110 51490 38162
rect 51886 38110 51938 38162
rect 53566 38110 53618 38162
rect 57710 38110 57762 38162
rect 14030 37998 14082 38050
rect 16606 37998 16658 38050
rect 17838 37998 17890 38050
rect 18734 37998 18786 38050
rect 20750 37998 20802 38050
rect 21870 37998 21922 38050
rect 23438 37998 23490 38050
rect 24782 37998 24834 38050
rect 25230 37998 25282 38050
rect 25454 37998 25506 38050
rect 26238 37998 26290 38050
rect 26574 37998 26626 38050
rect 27134 37998 27186 38050
rect 28590 37998 28642 38050
rect 29038 37998 29090 38050
rect 29262 37998 29314 38050
rect 29374 37998 29426 38050
rect 31166 37998 31218 38050
rect 31726 37998 31778 38050
rect 32062 37998 32114 38050
rect 32846 37998 32898 38050
rect 33070 37998 33122 38050
rect 34526 37998 34578 38050
rect 34862 37998 34914 38050
rect 35870 37998 35922 38050
rect 37550 37998 37602 38050
rect 37886 37998 37938 38050
rect 38110 37998 38162 38050
rect 42478 37998 42530 38050
rect 43262 37998 43314 38050
rect 43486 37998 43538 38050
rect 45390 37998 45442 38050
rect 51214 37998 51266 38050
rect 53454 37998 53506 38050
rect 54350 37998 54402 38050
rect 54574 37998 54626 38050
rect 55806 37998 55858 38050
rect 10222 37886 10274 37938
rect 18398 37886 18450 37938
rect 23998 37886 24050 37938
rect 28142 37886 28194 37938
rect 29710 37886 29762 37938
rect 34974 37886 35026 37938
rect 35646 37886 35698 37938
rect 42254 37886 42306 37938
rect 55246 37886 55298 37938
rect 10558 37774 10610 37826
rect 13470 37774 13522 37826
rect 15598 37774 15650 37826
rect 19742 37774 19794 37826
rect 20190 37774 20242 37826
rect 21310 37774 21362 37826
rect 25342 37774 25394 37826
rect 26014 37774 26066 37826
rect 26798 37774 26850 37826
rect 26910 37774 26962 37826
rect 27358 37774 27410 37826
rect 34302 37774 34354 37826
rect 37886 37774 37938 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 6974 37438 7026 37490
rect 7646 37438 7698 37490
rect 8654 37438 8706 37490
rect 15934 37438 15986 37490
rect 17614 37438 17666 37490
rect 18734 37438 18786 37490
rect 19070 37438 19122 37490
rect 22094 37438 22146 37490
rect 23550 37438 23602 37490
rect 23998 37438 24050 37490
rect 24334 37438 24386 37490
rect 27470 37438 27522 37490
rect 28254 37438 28306 37490
rect 33406 37438 33458 37490
rect 37662 37438 37714 37490
rect 40350 37438 40402 37490
rect 41358 37438 41410 37490
rect 50542 37438 50594 37490
rect 50654 37438 50706 37490
rect 54350 37438 54402 37490
rect 56030 37438 56082 37490
rect 1710 37326 1762 37378
rect 14030 37326 14082 37378
rect 15150 37326 15202 37378
rect 19630 37326 19682 37378
rect 24222 37326 24274 37378
rect 29710 37326 29762 37378
rect 30718 37326 30770 37378
rect 32174 37326 32226 37378
rect 33070 37326 33122 37378
rect 34078 37326 34130 37378
rect 37214 37326 37266 37378
rect 38446 37326 38498 37378
rect 39342 37326 39394 37378
rect 44270 37326 44322 37378
rect 49758 37326 49810 37378
rect 51662 37326 51714 37378
rect 54574 37326 54626 37378
rect 54798 37326 54850 37378
rect 55694 37326 55746 37378
rect 7198 37214 7250 37266
rect 8878 37214 8930 37266
rect 9662 37214 9714 37266
rect 10670 37214 10722 37266
rect 11118 37214 11170 37266
rect 13134 37214 13186 37266
rect 13582 37214 13634 37266
rect 15374 37214 15426 37266
rect 15598 37214 15650 37266
rect 18286 37214 18338 37266
rect 19854 37214 19906 37266
rect 20526 37214 20578 37266
rect 20750 37214 20802 37266
rect 21870 37214 21922 37266
rect 24558 37214 24610 37266
rect 26910 37214 26962 37266
rect 27246 37214 27298 37266
rect 27582 37214 27634 37266
rect 27806 37214 27858 37266
rect 28142 37214 28194 37266
rect 28478 37214 28530 37266
rect 28926 37214 28978 37266
rect 30046 37214 30098 37266
rect 30942 37214 30994 37266
rect 32062 37214 32114 37266
rect 33966 37214 34018 37266
rect 36206 37214 36258 37266
rect 38334 37214 38386 37266
rect 39006 37214 39058 37266
rect 39790 37214 39842 37266
rect 41022 37214 41074 37266
rect 41358 37214 41410 37266
rect 41694 37214 41746 37266
rect 42142 37214 42194 37266
rect 42366 37214 42418 37266
rect 44158 37214 44210 37266
rect 44494 37214 44546 37266
rect 44718 37214 44770 37266
rect 45278 37214 45330 37266
rect 45726 37214 45778 37266
rect 45950 37214 46002 37266
rect 50094 37214 50146 37266
rect 50766 37214 50818 37266
rect 51102 37214 51154 37266
rect 52894 37214 52946 37266
rect 54126 37214 54178 37266
rect 8206 37102 8258 37154
rect 9998 37102 10050 37154
rect 12686 37102 12738 37154
rect 17950 37102 18002 37154
rect 20190 37102 20242 37154
rect 29150 37102 29202 37154
rect 30158 37102 30210 37154
rect 31950 37102 32002 37154
rect 46062 37102 46114 37154
rect 49870 37102 49922 37154
rect 53006 37102 53058 37154
rect 2158 36990 2210 37042
rect 21198 36990 21250 37042
rect 40014 36990 40066 37042
rect 42030 36990 42082 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 13918 36654 13970 36706
rect 14590 36654 14642 36706
rect 22094 36654 22146 36706
rect 22318 36654 22370 36706
rect 26238 36654 26290 36706
rect 29486 36654 29538 36706
rect 35086 36654 35138 36706
rect 35422 36654 35474 36706
rect 36094 36654 36146 36706
rect 45950 36654 46002 36706
rect 50990 36654 51042 36706
rect 54238 36654 54290 36706
rect 1934 36542 1986 36594
rect 8990 36542 9042 36594
rect 11006 36542 11058 36594
rect 11790 36542 11842 36594
rect 18846 36542 18898 36594
rect 19406 36542 19458 36594
rect 20750 36542 20802 36594
rect 21534 36542 21586 36594
rect 23550 36542 23602 36594
rect 26574 36542 26626 36594
rect 29262 36542 29314 36594
rect 30382 36542 30434 36594
rect 31054 36542 31106 36594
rect 33518 36542 33570 36594
rect 41806 36542 41858 36594
rect 49310 36542 49362 36594
rect 51438 36542 51490 36594
rect 4286 36430 4338 36482
rect 8430 36430 8482 36482
rect 9438 36430 9490 36482
rect 9774 36430 9826 36482
rect 12126 36430 12178 36482
rect 12350 36430 12402 36482
rect 13470 36430 13522 36482
rect 13694 36430 13746 36482
rect 14142 36430 14194 36482
rect 15486 36430 15538 36482
rect 16382 36430 16434 36482
rect 17166 36430 17218 36482
rect 19742 36430 19794 36482
rect 20190 36430 20242 36482
rect 21870 36430 21922 36482
rect 22878 36430 22930 36482
rect 23998 36430 24050 36482
rect 24670 36430 24722 36482
rect 25566 36430 25618 36482
rect 27358 36430 27410 36482
rect 27582 36430 27634 36482
rect 27918 36430 27970 36482
rect 28254 36430 28306 36482
rect 29150 36430 29202 36482
rect 31390 36430 31442 36482
rect 32398 36430 32450 36482
rect 33294 36430 33346 36482
rect 33966 36430 34018 36482
rect 35198 36430 35250 36482
rect 35646 36430 35698 36482
rect 39342 36430 39394 36482
rect 41582 36430 41634 36482
rect 42254 36430 42306 36482
rect 44830 36430 44882 36482
rect 46062 36430 46114 36482
rect 47070 36430 47122 36482
rect 48526 36430 48578 36482
rect 49534 36430 49586 36482
rect 51214 36430 51266 36482
rect 53566 36430 53618 36482
rect 53902 36430 53954 36482
rect 55582 36430 55634 36482
rect 7534 36318 7586 36370
rect 12910 36318 12962 36370
rect 15374 36318 15426 36370
rect 15710 36318 15762 36370
rect 16158 36318 16210 36370
rect 18398 36318 18450 36370
rect 22766 36318 22818 36370
rect 24334 36318 24386 36370
rect 24894 36318 24946 36370
rect 26462 36318 26514 36370
rect 28142 36318 28194 36370
rect 30718 36318 30770 36370
rect 30942 36318 30994 36370
rect 32622 36318 32674 36370
rect 33182 36318 33234 36370
rect 34078 36318 34130 36370
rect 34414 36318 34466 36370
rect 35982 36318 36034 36370
rect 36094 36318 36146 36370
rect 37998 36318 38050 36370
rect 39118 36318 39170 36370
rect 42590 36318 42642 36370
rect 47294 36318 47346 36370
rect 49198 36318 49250 36370
rect 53790 36318 53842 36370
rect 54350 36318 54402 36370
rect 7870 36206 7922 36258
rect 17054 36206 17106 36258
rect 17726 36206 17778 36258
rect 18062 36206 18114 36258
rect 25678 36206 25730 36258
rect 27022 36206 27074 36258
rect 29934 36206 29986 36258
rect 34190 36206 34242 36258
rect 38110 36206 38162 36258
rect 38334 36206 38386 36258
rect 39566 36206 39618 36258
rect 56590 36206 56642 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 8206 35870 8258 35922
rect 14254 35870 14306 35922
rect 16270 35870 16322 35922
rect 17390 35870 17442 35922
rect 19070 35870 19122 35922
rect 19854 35870 19906 35922
rect 21422 35870 21474 35922
rect 24670 35870 24722 35922
rect 25342 35870 25394 35922
rect 27022 35870 27074 35922
rect 27246 35870 27298 35922
rect 28366 35870 28418 35922
rect 28814 35870 28866 35922
rect 29710 35870 29762 35922
rect 30158 35870 30210 35922
rect 34862 35870 34914 35922
rect 36766 35870 36818 35922
rect 41582 35870 41634 35922
rect 42366 35870 42418 35922
rect 10670 35758 10722 35810
rect 13582 35758 13634 35810
rect 14926 35758 14978 35810
rect 15710 35758 15762 35810
rect 22766 35758 22818 35810
rect 25230 35758 25282 35810
rect 26910 35758 26962 35810
rect 29486 35758 29538 35810
rect 30270 35758 30322 35810
rect 36206 35758 36258 35810
rect 37438 35758 37490 35810
rect 39454 35758 39506 35810
rect 41246 35758 41298 35810
rect 41358 35758 41410 35810
rect 43038 35758 43090 35810
rect 48078 35758 48130 35810
rect 49758 35758 49810 35810
rect 4286 35646 4338 35698
rect 6862 35646 6914 35698
rect 7422 35646 7474 35698
rect 8430 35646 8482 35698
rect 9998 35646 10050 35698
rect 11118 35646 11170 35698
rect 11678 35646 11730 35698
rect 12014 35646 12066 35698
rect 13246 35646 13298 35698
rect 14142 35646 14194 35698
rect 14814 35646 14866 35698
rect 15934 35646 15986 35698
rect 20414 35646 20466 35698
rect 25566 35646 25618 35698
rect 29374 35646 29426 35698
rect 29822 35646 29874 35698
rect 30382 35646 30434 35698
rect 33182 35646 33234 35698
rect 33630 35646 33682 35698
rect 34526 35646 34578 35698
rect 35310 35646 35362 35698
rect 35758 35646 35810 35698
rect 37214 35646 37266 35698
rect 37550 35646 37602 35698
rect 38334 35646 38386 35698
rect 38782 35646 38834 35698
rect 42814 35646 42866 35698
rect 45726 35646 45778 35698
rect 46286 35646 46338 35698
rect 47182 35646 47234 35698
rect 47406 35646 47458 35698
rect 49086 35646 49138 35698
rect 49534 35646 49586 35698
rect 52558 35646 52610 35698
rect 52782 35646 52834 35698
rect 53006 35646 53058 35698
rect 53230 35646 53282 35698
rect 53454 35646 53506 35698
rect 54238 35646 54290 35698
rect 55134 35646 55186 35698
rect 10110 35534 10162 35586
rect 12462 35534 12514 35586
rect 15374 35534 15426 35586
rect 17838 35534 17890 35586
rect 26014 35534 26066 35586
rect 32510 35534 32562 35586
rect 38670 35534 38722 35586
rect 43262 35534 43314 35586
rect 46734 35534 46786 35586
rect 52670 35534 52722 35586
rect 54350 35534 54402 35586
rect 1934 35422 1986 35474
rect 25678 35422 25730 35474
rect 26014 35422 26066 35474
rect 34302 35422 34354 35474
rect 36318 35422 36370 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 5518 35086 5570 35138
rect 20078 35086 20130 35138
rect 31278 35086 31330 35138
rect 33294 35086 33346 35138
rect 34078 35086 34130 35138
rect 44942 35086 44994 35138
rect 48862 35086 48914 35138
rect 12910 34974 12962 35026
rect 18062 34974 18114 35026
rect 18734 34974 18786 35026
rect 20750 34974 20802 35026
rect 22318 34974 22370 35026
rect 25902 34974 25954 35026
rect 27358 34974 27410 35026
rect 28702 34974 28754 35026
rect 30942 34974 30994 35026
rect 33854 34974 33906 35026
rect 38110 34974 38162 35026
rect 40574 34974 40626 35026
rect 50318 34974 50370 35026
rect 8654 34862 8706 34914
rect 8990 34862 9042 34914
rect 13470 34862 13522 34914
rect 14814 34862 14866 34914
rect 19406 34862 19458 34914
rect 19630 34862 19682 34914
rect 21870 34862 21922 34914
rect 22766 34862 22818 34914
rect 24222 34862 24274 34914
rect 24782 34862 24834 34914
rect 26350 34862 26402 34914
rect 27246 34862 27298 34914
rect 29150 34862 29202 34914
rect 30270 34862 30322 34914
rect 30494 34862 30546 34914
rect 31054 34862 31106 34914
rect 32286 34862 32338 34914
rect 37326 34862 37378 34914
rect 38222 34862 38274 34914
rect 39118 34862 39170 34914
rect 43374 34862 43426 34914
rect 44830 34862 44882 34914
rect 46846 34862 46898 34914
rect 47518 34862 47570 34914
rect 48078 34862 48130 34914
rect 48750 34862 48802 34914
rect 49198 34862 49250 34914
rect 49422 34862 49474 34914
rect 49758 34862 49810 34914
rect 52670 34862 52722 34914
rect 54686 34862 54738 34914
rect 9438 34750 9490 34802
rect 10446 34750 10498 34802
rect 13806 34750 13858 34802
rect 15038 34750 15090 34802
rect 18398 34750 18450 34802
rect 18622 34750 18674 34802
rect 26686 34750 26738 34802
rect 29486 34750 29538 34802
rect 32734 34750 32786 34802
rect 33518 34750 33570 34802
rect 37214 34750 37266 34802
rect 38558 34750 38610 34802
rect 44942 34750 44994 34802
rect 46510 34750 46562 34802
rect 49870 34750 49922 34802
rect 52782 34750 52834 34802
rect 55806 34750 55858 34802
rect 6302 34638 6354 34690
rect 9774 34638 9826 34690
rect 10110 34638 10162 34690
rect 10894 34638 10946 34690
rect 11342 34638 11394 34690
rect 14254 34638 14306 34690
rect 22990 34638 23042 34690
rect 32062 34638 32114 34690
rect 32846 34638 32898 34690
rect 34190 34638 34242 34690
rect 39454 34638 39506 34690
rect 43598 34638 43650 34690
rect 46622 34638 46674 34690
rect 52894 34638 52946 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 8318 34302 8370 34354
rect 9102 34302 9154 34354
rect 10558 34302 10610 34354
rect 11118 34302 11170 34354
rect 14478 34302 14530 34354
rect 16830 34302 16882 34354
rect 17390 34302 17442 34354
rect 21646 34302 21698 34354
rect 21758 34302 21810 34354
rect 22430 34302 22482 34354
rect 23214 34302 23266 34354
rect 23550 34302 23602 34354
rect 26014 34302 26066 34354
rect 26238 34302 26290 34354
rect 30158 34302 30210 34354
rect 30606 34302 30658 34354
rect 34190 34302 34242 34354
rect 35758 34302 35810 34354
rect 38894 34302 38946 34354
rect 43934 34302 43986 34354
rect 44494 34302 44546 34354
rect 46398 34302 46450 34354
rect 46510 34302 46562 34354
rect 47854 34302 47906 34354
rect 49870 34302 49922 34354
rect 50878 34302 50930 34354
rect 51998 34302 52050 34354
rect 53790 34302 53842 34354
rect 54350 34302 54402 34354
rect 54462 34302 54514 34354
rect 55582 34302 55634 34354
rect 18398 34190 18450 34242
rect 19070 34190 19122 34242
rect 19630 34190 19682 34242
rect 25678 34190 25730 34242
rect 29262 34190 29314 34242
rect 33630 34190 33682 34242
rect 34862 34190 34914 34242
rect 39230 34190 39282 34242
rect 40014 34190 40066 34242
rect 40350 34190 40402 34242
rect 45390 34190 45442 34242
rect 46846 34190 46898 34242
rect 46958 34190 47010 34242
rect 47630 34190 47682 34242
rect 50654 34190 50706 34242
rect 53006 34190 53058 34242
rect 54238 34190 54290 34242
rect 55246 34190 55298 34242
rect 5518 34078 5570 34130
rect 6078 34078 6130 34130
rect 9550 34078 9602 34130
rect 13694 34078 13746 34130
rect 14142 34078 14194 34130
rect 14702 34078 14754 34130
rect 17950 34078 18002 34130
rect 18734 34078 18786 34130
rect 19518 34078 19570 34130
rect 19742 34078 19794 34130
rect 19854 34078 19906 34130
rect 21086 34078 21138 34130
rect 21310 34078 21362 34130
rect 21534 34078 21586 34130
rect 25566 34078 25618 34130
rect 25902 34078 25954 34130
rect 26350 34078 26402 34130
rect 29710 34078 29762 34130
rect 30046 34078 30098 34130
rect 34750 34078 34802 34130
rect 36318 34078 36370 34130
rect 37886 34078 37938 34130
rect 38670 34078 38722 34130
rect 39454 34078 39506 34130
rect 41022 34078 41074 34130
rect 41358 34078 41410 34130
rect 45166 34078 45218 34130
rect 45950 34078 46002 34130
rect 46286 34078 46338 34130
rect 49646 34078 49698 34130
rect 50094 34078 50146 34130
rect 50206 34078 50258 34130
rect 50766 34078 50818 34130
rect 52446 34078 52498 34130
rect 9998 33966 10050 34018
rect 15262 33966 15314 34018
rect 31054 33966 31106 34018
rect 47966 33966 48018 34018
rect 51886 33966 51938 34018
rect 20190 33854 20242 33906
rect 20862 33854 20914 33906
rect 46958 33854 47010 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 14030 33518 14082 33570
rect 19518 33518 19570 33570
rect 24670 33518 24722 33570
rect 25230 33518 25282 33570
rect 26350 33518 26402 33570
rect 26462 33518 26514 33570
rect 37438 33518 37490 33570
rect 49310 33518 49362 33570
rect 51438 33518 51490 33570
rect 8318 33406 8370 33458
rect 18510 33406 18562 33458
rect 19294 33406 19346 33458
rect 21534 33406 21586 33458
rect 22990 33406 23042 33458
rect 23550 33406 23602 33458
rect 27582 33406 27634 33458
rect 45166 33406 45218 33458
rect 49982 33406 50034 33458
rect 50766 33406 50818 33458
rect 52782 33406 52834 33458
rect 57934 33406 57986 33458
rect 11678 33294 11730 33346
rect 12014 33294 12066 33346
rect 17166 33294 17218 33346
rect 17502 33294 17554 33346
rect 18846 33294 18898 33346
rect 19742 33294 19794 33346
rect 20078 33294 20130 33346
rect 21982 33294 22034 33346
rect 22654 33294 22706 33346
rect 24446 33294 24498 33346
rect 25006 33294 25058 33346
rect 25678 33294 25730 33346
rect 25902 33294 25954 33346
rect 26238 33294 26290 33346
rect 26686 33294 26738 33346
rect 36206 33294 36258 33346
rect 40462 33294 40514 33346
rect 40910 33294 40962 33346
rect 42478 33294 42530 33346
rect 43038 33294 43090 33346
rect 43710 33294 43762 33346
rect 45278 33294 45330 33346
rect 46510 33294 46562 33346
rect 47182 33294 47234 33346
rect 47518 33294 47570 33346
rect 48638 33294 48690 33346
rect 49534 33294 49586 33346
rect 53006 33294 53058 33346
rect 55582 33294 55634 33346
rect 1710 33182 1762 33234
rect 2046 33182 2098 33234
rect 8542 33182 8594 33234
rect 20414 33182 20466 33234
rect 22094 33182 22146 33234
rect 27022 33182 27074 33234
rect 36430 33182 36482 33234
rect 43150 33182 43202 33234
rect 48190 33182 48242 33234
rect 48526 33182 48578 33234
rect 49758 33182 49810 33234
rect 50094 33182 50146 33234
rect 50654 33182 50706 33234
rect 50878 33182 50930 33234
rect 51326 33182 51378 33234
rect 53678 33182 53730 33234
rect 54014 33182 54066 33234
rect 54350 33182 54402 33234
rect 2494 33070 2546 33122
rect 9102 33070 9154 33122
rect 12574 33070 12626 33122
rect 13582 33070 13634 33122
rect 14590 33070 14642 33122
rect 18958 33070 19010 33122
rect 19070 33070 19122 33122
rect 22206 33070 22258 33122
rect 23998 33070 24050 33122
rect 24334 33070 24386 33122
rect 26910 33070 26962 33122
rect 28590 33070 28642 33122
rect 29486 33070 29538 33122
rect 29822 33070 29874 33122
rect 30270 33070 30322 33122
rect 34302 33070 34354 33122
rect 37998 33070 38050 33122
rect 43486 33070 43538 33122
rect 47630 33070 47682 33122
rect 47854 33070 47906 33122
rect 48302 33070 48354 33122
rect 48974 33070 49026 33122
rect 49198 33070 49250 33122
rect 51438 33070 51490 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 19630 32734 19682 32786
rect 20526 32734 20578 32786
rect 22766 32734 22818 32786
rect 22990 32734 23042 32786
rect 24782 32734 24834 32786
rect 25454 32734 25506 32786
rect 29262 32734 29314 32786
rect 29822 32734 29874 32786
rect 36654 32734 36706 32786
rect 37214 32734 37266 32786
rect 43150 32734 43202 32786
rect 43710 32734 43762 32786
rect 47518 32734 47570 32786
rect 48078 32734 48130 32786
rect 50318 32734 50370 32786
rect 19854 32622 19906 32674
rect 23438 32622 23490 32674
rect 25230 32622 25282 32674
rect 37774 32622 37826 32674
rect 38110 32622 38162 32674
rect 38446 32622 38498 32674
rect 43598 32622 43650 32674
rect 43934 32622 43986 32674
rect 46958 32622 47010 32674
rect 47966 32622 48018 32674
rect 49646 32622 49698 32674
rect 16718 32510 16770 32562
rect 19966 32510 20018 32562
rect 22654 32510 22706 32562
rect 23102 32510 23154 32562
rect 25790 32510 25842 32562
rect 26126 32510 26178 32562
rect 26686 32510 26738 32562
rect 30158 32510 30210 32562
rect 33630 32510 33682 32562
rect 34078 32510 34130 32562
rect 37550 32510 37602 32562
rect 47182 32510 47234 32562
rect 48302 32510 48354 32562
rect 49758 32510 49810 32562
rect 49870 32510 49922 32562
rect 1822 32398 1874 32450
rect 11790 32398 11842 32450
rect 25566 32398 25618 32450
rect 30606 32398 30658 32450
rect 23550 32286 23602 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 48862 31950 48914 32002
rect 49198 31950 49250 32002
rect 37102 31838 37154 31890
rect 39006 31838 39058 31890
rect 39342 31838 39394 31890
rect 46174 31838 46226 31890
rect 48638 31838 48690 31890
rect 1822 31726 1874 31778
rect 24446 31726 24498 31778
rect 25006 31726 25058 31778
rect 30046 31726 30098 31778
rect 30494 31726 30546 31778
rect 33742 31726 33794 31778
rect 34190 31726 34242 31778
rect 34302 31726 34354 31778
rect 38670 31726 38722 31778
rect 2382 31614 2434 31666
rect 18510 31614 18562 31666
rect 19294 31614 19346 31666
rect 21310 31614 21362 31666
rect 32734 31614 32786 31666
rect 2046 31502 2098 31554
rect 4622 31502 4674 31554
rect 18174 31502 18226 31554
rect 18958 31502 19010 31554
rect 21982 31502 22034 31554
rect 25902 31502 25954 31554
rect 33518 31502 33570 31554
rect 34078 31502 34130 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 7870 31166 7922 31218
rect 8766 31166 8818 31218
rect 13022 31166 13074 31218
rect 16606 31166 16658 31218
rect 17502 31166 17554 31218
rect 25790 31166 25842 31218
rect 33742 31166 33794 31218
rect 38558 31166 38610 31218
rect 38782 31166 38834 31218
rect 39006 31166 39058 31218
rect 39678 31166 39730 31218
rect 41694 31166 41746 31218
rect 41918 31166 41970 31218
rect 45390 31166 45442 31218
rect 46174 31166 46226 31218
rect 9886 31054 9938 31106
rect 17838 31054 17890 31106
rect 21870 31054 21922 31106
rect 31838 31054 31890 31106
rect 40910 31054 40962 31106
rect 41246 31054 41298 31106
rect 47294 31054 47346 31106
rect 57822 31054 57874 31106
rect 4286 30942 4338 30994
rect 4846 30942 4898 30994
rect 5406 30942 5458 30994
rect 9662 30942 9714 30994
rect 15486 30942 15538 30994
rect 16158 30942 16210 30994
rect 18958 30942 19010 30994
rect 19406 30942 19458 30994
rect 25566 30942 25618 30994
rect 26910 30942 26962 30994
rect 33518 30942 33570 30994
rect 33854 30942 33906 30994
rect 41358 30942 41410 30994
rect 42030 30942 42082 30994
rect 42702 30942 42754 30994
rect 43038 30942 43090 30994
rect 46510 30942 46562 30994
rect 46734 30942 46786 30994
rect 58158 30942 58210 30994
rect 18622 30830 18674 30882
rect 26238 30830 26290 30882
rect 38670 30830 38722 30882
rect 39790 30830 39842 30882
rect 41022 30830 41074 30882
rect 57598 30830 57650 30882
rect 1934 30718 1986 30770
rect 8430 30718 8482 30770
rect 12462 30718 12514 30770
rect 39454 30718 39506 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 38894 30382 38946 30434
rect 42142 30382 42194 30434
rect 21758 30270 21810 30322
rect 23998 30270 24050 30322
rect 32062 30270 32114 30322
rect 4174 30158 4226 30210
rect 10782 30158 10834 30210
rect 11230 30158 11282 30210
rect 11790 30158 11842 30210
rect 13694 30158 13746 30210
rect 17614 30158 17666 30210
rect 17838 30158 17890 30210
rect 19182 30158 19234 30210
rect 19406 30158 19458 30210
rect 19630 30158 19682 30210
rect 20078 30158 20130 30210
rect 21982 30158 22034 30210
rect 23774 30158 23826 30210
rect 24222 30158 24274 30210
rect 25006 30158 25058 30210
rect 25342 30158 25394 30210
rect 32734 30158 32786 30210
rect 33966 30158 34018 30210
rect 38558 30158 38610 30210
rect 45950 30158 46002 30210
rect 2494 30046 2546 30098
rect 5630 30046 5682 30098
rect 5966 30046 6018 30098
rect 8542 30046 8594 30098
rect 13918 30046 13970 30098
rect 16942 30046 16994 30098
rect 18398 30046 18450 30098
rect 18510 30046 18562 30098
rect 21310 30046 21362 30098
rect 30718 30046 30770 30098
rect 31054 30046 31106 30098
rect 31726 30046 31778 30098
rect 32846 30046 32898 30098
rect 33294 30046 33346 30098
rect 40238 30046 40290 30098
rect 44158 30046 44210 30098
rect 44270 30046 44322 30098
rect 45614 30046 45666 30098
rect 45838 30046 45890 30098
rect 7758 29934 7810 29986
rect 18174 29934 18226 29986
rect 21534 29934 21586 29986
rect 21758 29934 21810 29986
rect 22542 29934 22594 29986
rect 24334 29934 24386 29986
rect 24446 29934 24498 29986
rect 27918 29934 27970 29986
rect 28478 29934 28530 29986
rect 33406 29934 33458 29986
rect 33630 29934 33682 29986
rect 37326 29934 37378 29986
rect 37662 29934 37714 29986
rect 39230 29934 39282 29986
rect 39566 29934 39618 29986
rect 43934 29934 43986 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 13694 29598 13746 29650
rect 19070 29598 19122 29650
rect 19966 29598 20018 29650
rect 21982 29598 22034 29650
rect 24670 29598 24722 29650
rect 25342 29598 25394 29650
rect 30830 29598 30882 29650
rect 31614 29598 31666 29650
rect 31726 29598 31778 29650
rect 36318 29598 36370 29650
rect 38446 29598 38498 29650
rect 46398 29598 46450 29650
rect 10110 29486 10162 29538
rect 14030 29486 14082 29538
rect 17950 29486 18002 29538
rect 19854 29486 19906 29538
rect 22206 29486 22258 29538
rect 22318 29486 22370 29538
rect 25230 29486 25282 29538
rect 26238 29486 26290 29538
rect 31950 29486 32002 29538
rect 32062 29486 32114 29538
rect 38334 29486 38386 29538
rect 38782 29486 38834 29538
rect 45614 29486 45666 29538
rect 4286 29374 4338 29426
rect 10558 29374 10610 29426
rect 11006 29374 11058 29426
rect 14366 29374 14418 29426
rect 15598 29374 15650 29426
rect 17614 29374 17666 29426
rect 17838 29374 17890 29426
rect 18174 29374 18226 29426
rect 18398 29374 18450 29426
rect 18846 29374 18898 29426
rect 21198 29374 21250 29426
rect 21646 29374 21698 29426
rect 25454 29374 25506 29426
rect 25678 29374 25730 29426
rect 28142 29374 28194 29426
rect 28590 29374 28642 29426
rect 33182 29374 33234 29426
rect 33742 29374 33794 29426
rect 39118 29374 39170 29426
rect 39454 29374 39506 29426
rect 42702 29374 42754 29426
rect 43262 29374 43314 29426
rect 9774 29262 9826 29314
rect 14926 29262 14978 29314
rect 16046 29262 16098 29314
rect 16718 29262 16770 29314
rect 18622 29262 18674 29314
rect 18958 29262 19010 29314
rect 19742 29262 19794 29314
rect 20750 29262 20802 29314
rect 22878 29262 22930 29314
rect 24222 29262 24274 29314
rect 37886 29262 37938 29314
rect 40238 29262 40290 29314
rect 1934 29150 1986 29202
rect 22318 29150 22370 29202
rect 24222 29150 24274 29202
rect 24446 29150 24498 29202
rect 24782 29150 24834 29202
rect 36878 29150 36930 29202
rect 39790 29150 39842 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 31390 28814 31442 28866
rect 1934 28702 1986 28754
rect 15038 28702 15090 28754
rect 18622 28702 18674 28754
rect 19294 28702 19346 28754
rect 21422 28702 21474 28754
rect 24222 28702 24274 28754
rect 25230 28702 25282 28754
rect 33070 28702 33122 28754
rect 33966 28702 34018 28754
rect 4286 28590 4338 28642
rect 6974 28590 7026 28642
rect 9774 28590 9826 28642
rect 10110 28590 10162 28642
rect 10558 28590 10610 28642
rect 12014 28590 12066 28642
rect 13470 28590 13522 28642
rect 13582 28590 13634 28642
rect 13918 28590 13970 28642
rect 14702 28590 14754 28642
rect 15486 28590 15538 28642
rect 16382 28590 16434 28642
rect 17838 28590 17890 28642
rect 19742 28590 19794 28642
rect 21310 28590 21362 28642
rect 21982 28590 22034 28642
rect 22318 28590 22370 28642
rect 22766 28590 22818 28642
rect 24558 28590 24610 28642
rect 25566 28590 25618 28642
rect 26126 28590 26178 28642
rect 29486 28590 29538 28642
rect 31054 28590 31106 28642
rect 31838 28590 31890 28642
rect 33518 28590 33570 28642
rect 37214 28590 37266 28642
rect 37326 28590 37378 28642
rect 37774 28590 37826 28642
rect 38222 28590 38274 28642
rect 11566 28478 11618 28530
rect 16046 28478 16098 28530
rect 16718 28478 16770 28530
rect 18174 28478 18226 28530
rect 20526 28478 20578 28530
rect 20638 28478 20690 28530
rect 24670 28478 24722 28530
rect 29150 28478 29202 28530
rect 32174 28478 32226 28530
rect 33182 28478 33234 28530
rect 37102 28478 37154 28530
rect 38558 28478 38610 28530
rect 7310 28366 7362 28418
rect 9214 28366 9266 28418
rect 13022 28366 13074 28418
rect 14254 28366 14306 28418
rect 17614 28366 17666 28418
rect 20302 28366 20354 28418
rect 20862 28366 20914 28418
rect 21534 28366 21586 28418
rect 28478 28366 28530 28418
rect 32958 28366 33010 28418
rect 58158 28366 58210 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 7310 28030 7362 28082
rect 8878 28030 8930 28082
rect 15598 28030 15650 28082
rect 18958 28030 19010 28082
rect 24670 28030 24722 28082
rect 26910 28030 26962 28082
rect 27694 28030 27746 28082
rect 29038 28030 29090 28082
rect 29822 28030 29874 28082
rect 30830 28030 30882 28082
rect 32622 28030 32674 28082
rect 35534 28030 35586 28082
rect 43934 28030 43986 28082
rect 8430 27918 8482 27970
rect 9550 27918 9602 27970
rect 9886 27918 9938 27970
rect 13246 27918 13298 27970
rect 13806 27918 13858 27970
rect 16270 27918 16322 27970
rect 26126 27918 26178 27970
rect 35646 27918 35698 27970
rect 36430 27918 36482 27970
rect 38222 27918 38274 27970
rect 38558 27918 38610 27970
rect 38670 27918 38722 27970
rect 4622 27806 4674 27858
rect 5070 27806 5122 27858
rect 10558 27806 10610 27858
rect 10782 27806 10834 27858
rect 11006 27806 11058 27858
rect 11230 27806 11282 27858
rect 12350 27806 12402 27858
rect 17390 27806 17442 27858
rect 23550 27806 23602 27858
rect 25678 27806 25730 27858
rect 28030 27806 28082 27858
rect 40798 27806 40850 27858
rect 41358 27806 41410 27858
rect 12126 27694 12178 27746
rect 14366 27694 14418 27746
rect 15150 27694 15202 27746
rect 16830 27694 16882 27746
rect 17950 27694 18002 27746
rect 18510 27694 18562 27746
rect 19518 27694 19570 27746
rect 19854 27694 19906 27746
rect 23998 27694 24050 27746
rect 25342 27694 25394 27746
rect 26462 27694 26514 27746
rect 28478 27694 28530 27746
rect 8094 27582 8146 27634
rect 8318 27582 8370 27634
rect 11678 27582 11730 27634
rect 12686 27582 12738 27634
rect 14030 27582 14082 27634
rect 35534 27582 35586 27634
rect 38558 27582 38610 27634
rect 44494 27582 44546 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 1934 27246 1986 27298
rect 11230 27246 11282 27298
rect 14254 27246 14306 27298
rect 16270 27246 16322 27298
rect 7646 27134 7698 27186
rect 8542 27134 8594 27186
rect 9550 27134 9602 27186
rect 14030 27134 14082 27186
rect 27694 27246 27746 27298
rect 16606 27134 16658 27186
rect 19854 27134 19906 27186
rect 21758 27134 21810 27186
rect 22318 27134 22370 27186
rect 22766 27134 22818 27186
rect 24222 27134 24274 27186
rect 27582 27134 27634 27186
rect 28478 27134 28530 27186
rect 29374 27134 29426 27186
rect 35758 27134 35810 27186
rect 37102 27134 37154 27186
rect 42590 27134 42642 27186
rect 4286 27022 4338 27074
rect 6638 27022 6690 27074
rect 7310 27022 7362 27074
rect 8206 27022 8258 27074
rect 10446 27022 10498 27074
rect 10670 27022 10722 27074
rect 10782 27022 10834 27074
rect 11566 27022 11618 27074
rect 12910 27022 12962 27074
rect 14030 27022 14082 27074
rect 14478 27022 14530 27074
rect 14926 27022 14978 27074
rect 15710 27022 15762 27074
rect 17166 27022 17218 27074
rect 17614 27022 17666 27074
rect 18062 27022 18114 27074
rect 18398 27022 18450 27074
rect 23214 27022 23266 27074
rect 25454 27022 25506 27074
rect 27246 27022 27298 27074
rect 28030 27022 28082 27074
rect 29150 27022 29202 27074
rect 30158 27022 30210 27074
rect 31278 27022 31330 27074
rect 31726 27022 31778 27074
rect 35198 27022 35250 27074
rect 36990 27022 37042 27074
rect 38782 27022 38834 27074
rect 39230 27022 39282 27074
rect 43038 27022 43090 27074
rect 43486 27022 43538 27074
rect 8990 26910 9042 26962
rect 12126 26910 12178 26962
rect 13470 26910 13522 26962
rect 13582 26910 13634 26962
rect 13694 26910 13746 26962
rect 16046 26910 16098 26962
rect 18846 26910 18898 26962
rect 20414 26910 20466 26962
rect 21310 26910 21362 26962
rect 23550 26910 23602 26962
rect 25790 26910 25842 26962
rect 27134 26910 27186 26962
rect 29262 26910 29314 26962
rect 30718 26910 30770 26962
rect 33966 26910 34018 26962
rect 34974 26910 35026 26962
rect 37438 26910 37490 26962
rect 41470 26910 41522 26962
rect 6862 26798 6914 26850
rect 19406 26798 19458 26850
rect 20750 26798 20802 26850
rect 34750 26798 34802 26850
rect 37214 26798 37266 26850
rect 42254 26798 42306 26850
rect 58158 26798 58210 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 1710 26462 1762 26514
rect 16270 26462 16322 26514
rect 39790 26462 39842 26514
rect 45166 26462 45218 26514
rect 5070 26350 5122 26402
rect 6078 26350 6130 26402
rect 15598 26350 15650 26402
rect 20526 26350 20578 26402
rect 24334 26350 24386 26402
rect 27694 26350 27746 26402
rect 39230 26350 39282 26402
rect 58158 26350 58210 26402
rect 4846 26238 4898 26290
rect 8094 26238 8146 26290
rect 10110 26238 10162 26290
rect 10334 26238 10386 26290
rect 12238 26238 12290 26290
rect 13806 26238 13858 26290
rect 14254 26238 14306 26290
rect 14702 26238 14754 26290
rect 15262 26238 15314 26290
rect 16158 26238 16210 26290
rect 18286 26238 18338 26290
rect 18622 26238 18674 26290
rect 19070 26238 19122 26290
rect 20190 26238 20242 26290
rect 21534 26238 21586 26290
rect 22206 26238 22258 26290
rect 22990 26238 23042 26290
rect 24446 26238 24498 26290
rect 26462 26238 26514 26290
rect 28254 26238 28306 26290
rect 29150 26238 29202 26290
rect 30382 26238 30434 26290
rect 31054 26238 31106 26290
rect 31278 26238 31330 26290
rect 38894 26238 38946 26290
rect 42254 26238 42306 26290
rect 42814 26238 42866 26290
rect 5966 26126 6018 26178
rect 6862 26126 6914 26178
rect 8654 26126 8706 26178
rect 9774 26126 9826 26178
rect 11678 26126 11730 26178
rect 12686 26126 12738 26178
rect 13470 26126 13522 26178
rect 16830 26126 16882 26178
rect 17838 26126 17890 26178
rect 19406 26126 19458 26178
rect 19742 26126 19794 26178
rect 20862 26126 20914 26178
rect 23774 26126 23826 26178
rect 26350 26126 26402 26178
rect 2158 26014 2210 26066
rect 13694 26014 13746 26066
rect 28478 26014 28530 26066
rect 31614 26014 31666 26066
rect 45950 26014 46002 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 7086 25678 7138 25730
rect 7422 25678 7474 25730
rect 9326 25678 9378 25730
rect 11342 25678 11394 25730
rect 30494 25678 30546 25730
rect 31278 25678 31330 25730
rect 42814 25678 42866 25730
rect 11902 25566 11954 25618
rect 15374 25566 15426 25618
rect 16494 25566 16546 25618
rect 17390 25566 17442 25618
rect 21758 25566 21810 25618
rect 22766 25566 22818 25618
rect 25902 25566 25954 25618
rect 28142 25566 28194 25618
rect 30718 25566 30770 25618
rect 31278 25566 31330 25618
rect 31614 25566 31666 25618
rect 32174 25566 32226 25618
rect 36094 25566 36146 25618
rect 42366 25566 42418 25618
rect 57934 25566 57986 25618
rect 5966 25454 6018 25506
rect 9438 25454 9490 25506
rect 9886 25454 9938 25506
rect 10670 25454 10722 25506
rect 11006 25454 11058 25506
rect 12238 25454 12290 25506
rect 12686 25454 12738 25506
rect 13918 25454 13970 25506
rect 14142 25454 14194 25506
rect 15262 25454 15314 25506
rect 15934 25454 15986 25506
rect 17054 25454 17106 25506
rect 17950 25454 18002 25506
rect 20190 25454 20242 25506
rect 22318 25454 22370 25506
rect 23214 25454 23266 25506
rect 23886 25454 23938 25506
rect 25118 25454 25170 25506
rect 26126 25454 26178 25506
rect 28590 25454 28642 25506
rect 29150 25454 29202 25506
rect 30046 25454 30098 25506
rect 31838 25454 31890 25506
rect 34414 25454 34466 25506
rect 35086 25454 35138 25506
rect 35534 25454 35586 25506
rect 37998 25454 38050 25506
rect 38558 25454 38610 25506
rect 43934 25454 43986 25506
rect 46846 25454 46898 25506
rect 55582 25454 55634 25506
rect 5630 25342 5682 25394
rect 6862 25342 6914 25394
rect 9326 25342 9378 25394
rect 10334 25342 10386 25394
rect 12462 25342 12514 25394
rect 12910 25342 12962 25394
rect 13022 25342 13074 25394
rect 15486 25342 15538 25394
rect 16270 25342 16322 25394
rect 17614 25342 17666 25394
rect 17726 25342 17778 25394
rect 19294 25342 19346 25394
rect 21534 25342 21586 25394
rect 29262 25342 29314 25394
rect 35758 25342 35810 25394
rect 37326 25342 37378 25394
rect 38670 25342 38722 25394
rect 42814 25342 42866 25394
rect 42926 25342 42978 25394
rect 43150 25342 43202 25394
rect 43374 25342 43426 25394
rect 43486 25342 43538 25394
rect 47070 25342 47122 25394
rect 8990 25230 9042 25282
rect 13582 25230 13634 25282
rect 18398 25230 18450 25282
rect 18958 25230 19010 25282
rect 24558 25230 24610 25282
rect 30158 25230 30210 25282
rect 34078 25230 34130 25282
rect 36206 25230 36258 25282
rect 36990 25230 37042 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 7422 24894 7474 24946
rect 16158 24894 16210 24946
rect 17502 24894 17554 24946
rect 24670 24894 24722 24946
rect 27470 24894 27522 24946
rect 27806 24894 27858 24946
rect 29262 24894 29314 24946
rect 29710 24894 29762 24946
rect 30606 24894 30658 24946
rect 38894 24894 38946 24946
rect 8990 24782 9042 24834
rect 12014 24782 12066 24834
rect 12686 24782 12738 24834
rect 13022 24782 13074 24834
rect 14926 24782 14978 24834
rect 20974 24782 21026 24834
rect 23438 24782 23490 24834
rect 24110 24782 24162 24834
rect 28366 24782 28418 24834
rect 28702 24782 28754 24834
rect 33406 24782 33458 24834
rect 36094 24782 36146 24834
rect 38782 24782 38834 24834
rect 41358 24782 41410 24834
rect 43262 24782 43314 24834
rect 46846 24782 46898 24834
rect 6078 24670 6130 24722
rect 8542 24670 8594 24722
rect 9550 24670 9602 24722
rect 10110 24670 10162 24722
rect 12910 24670 12962 24722
rect 13470 24670 13522 24722
rect 15822 24670 15874 24722
rect 17838 24670 17890 24722
rect 18398 24670 18450 24722
rect 20190 24670 20242 24722
rect 21870 24670 21922 24722
rect 22430 24670 22482 24722
rect 23214 24670 23266 24722
rect 25566 24670 25618 24722
rect 26574 24670 26626 24722
rect 30942 24670 30994 24722
rect 31166 24670 31218 24722
rect 31838 24670 31890 24722
rect 33182 24670 33234 24722
rect 34974 24670 35026 24722
rect 35534 24670 35586 24722
rect 36878 24670 36930 24722
rect 37886 24670 37938 24722
rect 38110 24670 38162 24722
rect 39118 24670 39170 24722
rect 42254 24670 42306 24722
rect 42702 24670 42754 24722
rect 46174 24670 46226 24722
rect 46622 24670 46674 24722
rect 6638 24558 6690 24610
rect 7870 24558 7922 24610
rect 11006 24558 11058 24610
rect 14366 24558 14418 24610
rect 16606 24558 16658 24610
rect 21198 24558 21250 24610
rect 23326 24558 23378 24610
rect 26014 24558 26066 24610
rect 26910 24558 26962 24610
rect 30158 24558 30210 24610
rect 35982 24558 36034 24610
rect 37326 24558 37378 24610
rect 41694 24558 41746 24610
rect 42814 24558 42866 24610
rect 43374 24558 43426 24610
rect 1710 24446 1762 24498
rect 26462 24446 26514 24498
rect 31390 24446 31442 24498
rect 38446 24446 38498 24498
rect 43486 24446 43538 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 5742 24110 5794 24162
rect 19406 24110 19458 24162
rect 46622 24110 46674 24162
rect 46958 24110 47010 24162
rect 47518 24110 47570 24162
rect 5630 23998 5682 24050
rect 6414 23998 6466 24050
rect 18510 23998 18562 24050
rect 19294 23998 19346 24050
rect 20750 23998 20802 24050
rect 28142 23998 28194 24050
rect 31166 23998 31218 24050
rect 40798 23998 40850 24050
rect 43486 23998 43538 24050
rect 45838 23998 45890 24050
rect 46398 23998 46450 24050
rect 57934 23998 57986 24050
rect 7310 23886 7362 23938
rect 8430 23886 8482 23938
rect 9326 23886 9378 23938
rect 9662 23886 9714 23938
rect 11006 23886 11058 23938
rect 11902 23886 11954 23938
rect 14478 23886 14530 23938
rect 14814 23886 14866 23938
rect 15374 23886 15426 23938
rect 15934 23886 15986 23938
rect 16942 23886 16994 23938
rect 17838 23886 17890 23938
rect 18398 23886 18450 23938
rect 19406 23886 19458 23938
rect 22094 23886 22146 23938
rect 22542 23886 22594 23938
rect 22990 23886 23042 23938
rect 24446 23886 24498 23938
rect 26350 23886 26402 23938
rect 27470 23886 27522 23938
rect 28478 23886 28530 23938
rect 29150 23886 29202 23938
rect 29598 23886 29650 23938
rect 31390 23886 31442 23938
rect 33406 23886 33458 23938
rect 41134 23886 41186 23938
rect 41694 23886 41746 23938
rect 42030 23886 42082 23938
rect 42590 23886 42642 23938
rect 43374 23886 43426 23938
rect 47294 23886 47346 23938
rect 55582 23886 55634 23938
rect 9998 23774 10050 23826
rect 11342 23774 11394 23826
rect 12910 23774 12962 23826
rect 15710 23774 15762 23826
rect 16830 23774 16882 23826
rect 23998 23774 24050 23826
rect 26126 23774 26178 23826
rect 31502 23774 31554 23826
rect 34526 23774 34578 23826
rect 44270 23774 44322 23826
rect 45950 23774 46002 23826
rect 50094 23774 50146 23826
rect 13918 23662 13970 23714
rect 17726 23662 17778 23714
rect 21310 23662 21362 23714
rect 25454 23662 25506 23714
rect 27134 23662 27186 23714
rect 35086 23662 35138 23714
rect 40686 23662 40738 23714
rect 42366 23662 42418 23714
rect 42478 23662 42530 23714
rect 45502 23662 45554 23714
rect 45726 23662 45778 23714
rect 47854 23662 47906 23714
rect 49758 23662 49810 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 17614 23326 17666 23378
rect 21870 23326 21922 23378
rect 40910 23326 40962 23378
rect 42590 23326 42642 23378
rect 43150 23326 43202 23378
rect 7758 23214 7810 23266
rect 11678 23214 11730 23266
rect 18846 23214 18898 23266
rect 22430 23214 22482 23266
rect 22654 23214 22706 23266
rect 24670 23214 24722 23266
rect 26014 23214 26066 23266
rect 26350 23214 26402 23266
rect 29486 23214 29538 23266
rect 31390 23214 31442 23266
rect 33742 23214 33794 23266
rect 41246 23214 41298 23266
rect 42814 23214 42866 23266
rect 44942 23214 44994 23266
rect 49758 23214 49810 23266
rect 5070 23102 5122 23154
rect 5630 23102 5682 23154
rect 8430 23102 8482 23154
rect 10222 23102 10274 23154
rect 11006 23102 11058 23154
rect 12798 23102 12850 23154
rect 14142 23102 14194 23154
rect 14926 23102 14978 23154
rect 18062 23102 18114 23154
rect 19630 23102 19682 23154
rect 20638 23102 20690 23154
rect 21422 23102 21474 23154
rect 23102 23102 23154 23154
rect 24334 23102 24386 23154
rect 25678 23102 25730 23154
rect 26686 23102 26738 23154
rect 27470 23102 27522 23154
rect 28254 23102 28306 23154
rect 29934 23102 29986 23154
rect 30942 23102 30994 23154
rect 31278 23102 31330 23154
rect 31950 23102 32002 23154
rect 32510 23102 32562 23154
rect 33518 23102 33570 23154
rect 33630 23102 33682 23154
rect 35086 23102 35138 23154
rect 35758 23102 35810 23154
rect 38894 23102 38946 23154
rect 41918 23102 41970 23154
rect 42142 23102 42194 23154
rect 45390 23102 45442 23154
rect 46174 23102 46226 23154
rect 49086 23102 49138 23154
rect 6526 22990 6578 23042
rect 7198 22990 7250 23042
rect 7758 22990 7810 23042
rect 9998 22990 10050 23042
rect 10894 22990 10946 23042
rect 12238 22990 12290 23042
rect 15710 22990 15762 23042
rect 16158 22990 16210 23042
rect 16606 22990 16658 23042
rect 22766 22990 22818 23042
rect 24446 22990 24498 23042
rect 25342 22990 25394 23042
rect 26910 22990 26962 23042
rect 29038 22990 29090 23042
rect 34302 22990 34354 23042
rect 34862 22990 34914 23042
rect 38334 22990 38386 23042
rect 39118 22990 39170 23042
rect 41694 22990 41746 23042
rect 44606 22990 44658 23042
rect 46398 22990 46450 23042
rect 46846 22990 46898 23042
rect 48862 22990 48914 23042
rect 13918 22878 13970 22930
rect 15486 22878 15538 22930
rect 16382 22878 16434 22930
rect 23326 22878 23378 22930
rect 23662 22878 23714 22930
rect 33070 22878 33122 22930
rect 39342 22878 39394 22930
rect 45054 22878 45106 22930
rect 45502 22878 45554 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 26574 22542 26626 22594
rect 29150 22542 29202 22594
rect 10110 22430 10162 22482
rect 16718 22430 16770 22482
rect 17614 22430 17666 22482
rect 20302 22430 20354 22482
rect 20750 22430 20802 22482
rect 25454 22430 25506 22482
rect 45614 22542 45666 22594
rect 49198 22542 49250 22594
rect 29822 22430 29874 22482
rect 31502 22430 31554 22482
rect 33406 22430 33458 22482
rect 35198 22430 35250 22482
rect 36206 22430 36258 22482
rect 37774 22430 37826 22482
rect 38334 22430 38386 22482
rect 39230 22430 39282 22482
rect 40462 22430 40514 22482
rect 48974 22430 49026 22482
rect 57934 22430 57986 22482
rect 6078 22318 6130 22370
rect 6638 22318 6690 22370
rect 6974 22318 7026 22370
rect 8542 22318 8594 22370
rect 8990 22318 9042 22370
rect 10558 22318 10610 22370
rect 12462 22318 12514 22370
rect 14142 22318 14194 22370
rect 15822 22318 15874 22370
rect 16270 22318 16322 22370
rect 17278 22318 17330 22370
rect 18062 22318 18114 22370
rect 19182 22318 19234 22370
rect 19742 22318 19794 22370
rect 20190 22318 20242 22370
rect 21422 22318 21474 22370
rect 21646 22318 21698 22370
rect 23550 22318 23602 22370
rect 25902 22318 25954 22370
rect 26126 22318 26178 22370
rect 26462 22318 26514 22370
rect 26686 22318 26738 22370
rect 27022 22318 27074 22370
rect 27582 22318 27634 22370
rect 28478 22318 28530 22370
rect 29822 22318 29874 22370
rect 31950 22318 32002 22370
rect 33854 22318 33906 22370
rect 34974 22318 35026 22370
rect 35758 22318 35810 22370
rect 35982 22318 36034 22370
rect 39006 22318 39058 22370
rect 40014 22318 40066 22370
rect 44942 22318 44994 22370
rect 45278 22318 45330 22370
rect 45726 22318 45778 22370
rect 46398 22318 46450 22370
rect 55582 22318 55634 22370
rect 7534 22206 7586 22258
rect 11566 22206 11618 22258
rect 12014 22206 12066 22258
rect 13470 22206 13522 22258
rect 18174 22206 18226 22258
rect 24670 22206 24722 22258
rect 28030 22206 28082 22258
rect 29262 22206 29314 22258
rect 30942 22206 30994 22258
rect 32398 22206 32450 22258
rect 37214 22206 37266 22258
rect 37326 22206 37378 22258
rect 37438 22206 37490 22258
rect 39678 22206 39730 22258
rect 46174 22206 46226 22258
rect 8094 22094 8146 22146
rect 8318 22094 8370 22146
rect 9326 22094 9378 22146
rect 15710 22094 15762 22146
rect 18958 22094 19010 22146
rect 24894 22094 24946 22146
rect 36990 22094 37042 22146
rect 45502 22094 45554 22146
rect 46286 22094 46338 22146
rect 49534 22094 49586 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 5630 21758 5682 21810
rect 5854 21758 5906 21810
rect 10334 21758 10386 21810
rect 17726 21758 17778 21810
rect 22430 21758 22482 21810
rect 26014 21758 26066 21810
rect 26798 21758 26850 21810
rect 27806 21758 27858 21810
rect 28366 21758 28418 21810
rect 29598 21758 29650 21810
rect 32062 21758 32114 21810
rect 33854 21758 33906 21810
rect 35198 21758 35250 21810
rect 41694 21758 41746 21810
rect 42142 21758 42194 21810
rect 42478 21758 42530 21810
rect 51102 21758 51154 21810
rect 58158 21758 58210 21810
rect 1710 21646 1762 21698
rect 11566 21646 11618 21698
rect 14254 21646 14306 21698
rect 20190 21646 20242 21698
rect 21198 21646 21250 21698
rect 26238 21646 26290 21698
rect 28926 21646 28978 21698
rect 29150 21646 29202 21698
rect 31054 21646 31106 21698
rect 31166 21646 31218 21698
rect 32398 21646 32450 21698
rect 35086 21646 35138 21698
rect 37550 21646 37602 21698
rect 42814 21646 42866 21698
rect 43038 21646 43090 21698
rect 43374 21646 43426 21698
rect 6414 21534 6466 21586
rect 7310 21534 7362 21586
rect 11230 21534 11282 21586
rect 14814 21534 14866 21586
rect 16158 21534 16210 21586
rect 18622 21534 18674 21586
rect 19070 21534 19122 21586
rect 20302 21534 20354 21586
rect 21086 21534 21138 21586
rect 21870 21534 21922 21586
rect 23102 21534 23154 21586
rect 23438 21534 23490 21586
rect 24334 21534 24386 21586
rect 25230 21534 25282 21586
rect 25342 21534 25394 21586
rect 25454 21534 25506 21586
rect 25790 21534 25842 21586
rect 26350 21534 26402 21586
rect 28590 21534 28642 21586
rect 30046 21534 30098 21586
rect 30830 21534 30882 21586
rect 33070 21534 33122 21586
rect 33294 21534 33346 21586
rect 33518 21534 33570 21586
rect 33742 21534 33794 21586
rect 34078 21534 34130 21586
rect 34974 21534 35026 21586
rect 38670 21534 38722 21586
rect 39566 21534 39618 21586
rect 41582 21534 41634 21586
rect 49758 21534 49810 21586
rect 50430 21534 50482 21586
rect 50766 21534 50818 21586
rect 6974 21422 7026 21474
rect 7982 21422 8034 21474
rect 8990 21422 9042 21474
rect 10110 21422 10162 21474
rect 10894 21422 10946 21474
rect 11902 21422 11954 21474
rect 12462 21422 12514 21474
rect 12910 21422 12962 21474
rect 15038 21422 15090 21474
rect 15598 21422 15650 21474
rect 16606 21422 16658 21474
rect 18286 21422 18338 21474
rect 19854 21422 19906 21474
rect 23886 21422 23938 21474
rect 27246 21422 27298 21474
rect 30606 21422 30658 21474
rect 31726 21422 31778 21474
rect 34638 21422 34690 21474
rect 39230 21422 39282 21474
rect 43262 21422 43314 21474
rect 49534 21422 49586 21474
rect 24222 21310 24274 21362
rect 32510 21310 32562 21362
rect 41694 21310 41746 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 17054 20974 17106 21026
rect 31838 20974 31890 21026
rect 33854 20974 33906 21026
rect 35646 20974 35698 21026
rect 6974 20862 7026 20914
rect 8990 20862 9042 20914
rect 11342 20862 11394 20914
rect 12238 20862 12290 20914
rect 13918 20862 13970 20914
rect 16718 20862 16770 20914
rect 18174 20862 18226 20914
rect 35870 20862 35922 20914
rect 36206 20862 36258 20914
rect 37662 20862 37714 20914
rect 38670 20862 38722 20914
rect 42366 20862 42418 20914
rect 43710 20862 43762 20914
rect 44046 20862 44098 20914
rect 48638 20862 48690 20914
rect 49534 20862 49586 20914
rect 7534 20750 7586 20802
rect 8094 20750 8146 20802
rect 10222 20750 10274 20802
rect 11790 20750 11842 20802
rect 13694 20750 13746 20802
rect 15822 20750 15874 20802
rect 16270 20750 16322 20802
rect 16494 20750 16546 20802
rect 17390 20750 17442 20802
rect 17614 20750 17666 20802
rect 19406 20750 19458 20802
rect 22206 20750 22258 20802
rect 23774 20750 23826 20802
rect 25342 20750 25394 20802
rect 26238 20750 26290 20802
rect 27246 20750 27298 20802
rect 28030 20750 28082 20802
rect 28478 20750 28530 20802
rect 29598 20750 29650 20802
rect 30718 20750 30770 20802
rect 31614 20750 31666 20802
rect 33518 20750 33570 20802
rect 34638 20750 34690 20802
rect 35086 20750 35138 20802
rect 36318 20750 36370 20802
rect 38110 20750 38162 20802
rect 39678 20750 39730 20802
rect 41134 20750 41186 20802
rect 41358 20750 41410 20802
rect 41582 20750 41634 20802
rect 41694 20750 41746 20802
rect 42814 20750 42866 20802
rect 43262 20750 43314 20802
rect 47294 20750 47346 20802
rect 47966 20750 48018 20802
rect 48862 20750 48914 20802
rect 49758 20750 49810 20802
rect 6302 20638 6354 20690
rect 8654 20638 8706 20690
rect 12686 20638 12738 20690
rect 13470 20638 13522 20690
rect 16830 20638 16882 20690
rect 19294 20638 19346 20690
rect 22318 20638 22370 20690
rect 26014 20638 26066 20690
rect 26798 20638 26850 20690
rect 27022 20638 27074 20690
rect 31950 20638 32002 20690
rect 34974 20638 35026 20690
rect 39902 20638 39954 20690
rect 40350 20638 40402 20690
rect 40910 20638 40962 20690
rect 45614 20638 45666 20690
rect 46062 20638 46114 20690
rect 46174 20638 46226 20690
rect 46734 20638 46786 20690
rect 50318 20638 50370 20690
rect 9550 20526 9602 20578
rect 12798 20526 12850 20578
rect 13022 20526 13074 20578
rect 18622 20526 18674 20578
rect 20638 20526 20690 20578
rect 21646 20526 21698 20578
rect 22430 20526 22482 20578
rect 36094 20526 36146 20578
rect 41918 20526 41970 20578
rect 44158 20526 44210 20578
rect 45838 20526 45890 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 16606 20190 16658 20242
rect 18958 20190 19010 20242
rect 22094 20190 22146 20242
rect 23326 20190 23378 20242
rect 30718 20190 30770 20242
rect 31726 20190 31778 20242
rect 31838 20190 31890 20242
rect 34862 20190 34914 20242
rect 40238 20190 40290 20242
rect 58158 20190 58210 20242
rect 5294 20078 5346 20130
rect 9774 20078 9826 20130
rect 15150 20078 15202 20130
rect 18062 20078 18114 20130
rect 19182 20078 19234 20130
rect 19742 20078 19794 20130
rect 22430 20078 22482 20130
rect 24222 20078 24274 20130
rect 25566 20078 25618 20130
rect 26574 20078 26626 20130
rect 27470 20078 27522 20130
rect 28142 20078 28194 20130
rect 28590 20078 28642 20130
rect 33294 20078 33346 20130
rect 33630 20078 33682 20130
rect 34526 20078 34578 20130
rect 36206 20078 36258 20130
rect 39454 20078 39506 20130
rect 41582 20078 41634 20130
rect 46174 20078 46226 20130
rect 46734 20078 46786 20130
rect 49198 20078 49250 20130
rect 49310 20078 49362 20130
rect 5854 19966 5906 20018
rect 7086 19966 7138 20018
rect 8542 19966 8594 20018
rect 9550 19966 9602 20018
rect 10894 19966 10946 20018
rect 12462 19966 12514 20018
rect 13022 19966 13074 20018
rect 13470 19966 13522 20018
rect 13694 19966 13746 20018
rect 16606 19966 16658 20018
rect 18622 19966 18674 20018
rect 19406 19966 19458 20018
rect 20078 19966 20130 20018
rect 21086 19966 21138 20018
rect 21310 19966 21362 20018
rect 22318 19966 22370 20018
rect 23438 19966 23490 20018
rect 23998 19966 24050 20018
rect 24446 19966 24498 20018
rect 24558 19966 24610 20018
rect 25342 19966 25394 20018
rect 26238 19966 26290 20018
rect 27582 19966 27634 20018
rect 27694 19966 27746 20018
rect 28814 19966 28866 20018
rect 30830 19966 30882 20018
rect 31614 19966 31666 20018
rect 31950 19966 32002 20018
rect 32174 19966 32226 20018
rect 33070 19966 33122 20018
rect 35982 19966 36034 20018
rect 36542 19966 36594 20018
rect 37886 19966 37938 20018
rect 38334 19966 38386 20018
rect 38558 19966 38610 20018
rect 39342 19966 39394 20018
rect 40126 19966 40178 20018
rect 41918 19966 41970 20018
rect 42702 19966 42754 20018
rect 42926 19966 42978 20018
rect 44718 19966 44770 20018
rect 44942 19966 44994 20018
rect 46062 19966 46114 20018
rect 46846 19966 46898 20018
rect 47518 19966 47570 20018
rect 47966 19966 48018 20018
rect 49534 19966 49586 20018
rect 4958 19854 5010 19906
rect 7422 19854 7474 19906
rect 7646 19854 7698 19906
rect 8430 19854 8482 19906
rect 10222 19854 10274 19906
rect 11342 19854 11394 19906
rect 17614 19854 17666 19906
rect 20414 19854 20466 19906
rect 20862 19854 20914 19906
rect 26014 19854 26066 19906
rect 34302 19854 34354 19906
rect 37102 19854 37154 19906
rect 38446 19854 38498 19906
rect 45950 19854 46002 19906
rect 8766 19742 8818 19794
rect 18958 19742 19010 19794
rect 43710 19742 43762 19794
rect 47070 19742 47122 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 6750 19406 6802 19458
rect 17502 19406 17554 19458
rect 17838 19406 17890 19458
rect 23886 19406 23938 19458
rect 23998 19406 24050 19458
rect 24222 19406 24274 19458
rect 40686 19406 40738 19458
rect 43710 19406 43762 19458
rect 44270 19406 44322 19458
rect 46958 19406 47010 19458
rect 49198 19406 49250 19458
rect 11566 19294 11618 19346
rect 13582 19294 13634 19346
rect 14142 19294 14194 19346
rect 15038 19294 15090 19346
rect 18398 19294 18450 19346
rect 21422 19294 21474 19346
rect 25118 19294 25170 19346
rect 27582 19294 27634 19346
rect 28142 19294 28194 19346
rect 32734 19294 32786 19346
rect 38222 19294 38274 19346
rect 44046 19294 44098 19346
rect 48974 19294 49026 19346
rect 50094 19294 50146 19346
rect 5630 19182 5682 19234
rect 6526 19182 6578 19234
rect 7646 19182 7698 19234
rect 7870 19182 7922 19234
rect 8318 19182 8370 19234
rect 9102 19182 9154 19234
rect 9662 19182 9714 19234
rect 11454 19182 11506 19234
rect 12014 19182 12066 19234
rect 14254 19182 14306 19234
rect 15262 19182 15314 19234
rect 15934 19182 15986 19234
rect 18734 19182 18786 19234
rect 19182 19182 19234 19234
rect 20302 19182 20354 19234
rect 21870 19182 21922 19234
rect 22766 19182 22818 19234
rect 22990 19182 23042 19234
rect 25678 19182 25730 19234
rect 26014 19182 26066 19234
rect 26238 19182 26290 19234
rect 29262 19182 29314 19234
rect 29598 19182 29650 19234
rect 29934 19182 29986 19234
rect 36430 19182 36482 19234
rect 37438 19182 37490 19234
rect 38334 19182 38386 19234
rect 40014 19182 40066 19234
rect 43486 19182 43538 19234
rect 46286 19182 46338 19234
rect 46622 19182 46674 19234
rect 51438 19182 51490 19234
rect 7086 19070 7138 19122
rect 10894 19070 10946 19122
rect 15710 19070 15762 19122
rect 16270 19070 16322 19122
rect 16942 19070 16994 19122
rect 17278 19070 17330 19122
rect 19966 19070 20018 19122
rect 22318 19070 22370 19122
rect 22878 19070 22930 19122
rect 25902 19070 25954 19122
rect 37214 19070 37266 19122
rect 38558 19070 38610 19122
rect 40126 19070 40178 19122
rect 40238 19070 40290 19122
rect 44046 19070 44098 19122
rect 49534 19070 49586 19122
rect 50206 19070 50258 19122
rect 52110 19070 52162 19122
rect 52670 19070 52722 19122
rect 5966 18958 6018 19010
rect 7758 18958 7810 19010
rect 8990 18958 9042 19010
rect 9550 18958 9602 19010
rect 9774 18958 9826 19010
rect 18846 18958 18898 19010
rect 20414 18958 20466 19010
rect 23438 18958 23490 19010
rect 23886 18958 23938 19010
rect 25006 18958 25058 19010
rect 25230 18958 25282 19010
rect 27134 18958 27186 19010
rect 28590 18958 28642 19010
rect 29598 18958 29650 19010
rect 30382 18958 30434 19010
rect 31166 18958 31218 19010
rect 31614 18958 31666 19010
rect 33630 18958 33682 19010
rect 33966 18958 34018 19010
rect 35870 18958 35922 19010
rect 42366 18958 42418 19010
rect 46846 18958 46898 19010
rect 53006 18958 53058 19010
rect 58158 18958 58210 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 7310 18622 7362 18674
rect 11342 18622 11394 18674
rect 19406 18622 19458 18674
rect 24222 18622 24274 18674
rect 24446 18622 24498 18674
rect 24670 18622 24722 18674
rect 26686 18622 26738 18674
rect 28478 18622 28530 18674
rect 43598 18622 43650 18674
rect 5182 18510 5234 18562
rect 7198 18510 7250 18562
rect 7982 18510 8034 18562
rect 8318 18510 8370 18562
rect 8990 18510 9042 18562
rect 10334 18510 10386 18562
rect 15822 18510 15874 18562
rect 16270 18510 16322 18562
rect 16718 18510 16770 18562
rect 17614 18510 17666 18562
rect 18622 18510 18674 18562
rect 29486 18510 29538 18562
rect 30494 18510 30546 18562
rect 37550 18510 37602 18562
rect 43822 18510 43874 18562
rect 44046 18510 44098 18562
rect 49758 18510 49810 18562
rect 6078 18398 6130 18450
rect 6862 18398 6914 18450
rect 7534 18398 7586 18450
rect 7870 18398 7922 18450
rect 10446 18398 10498 18450
rect 13358 18398 13410 18450
rect 13694 18398 13746 18450
rect 14590 18398 14642 18450
rect 15486 18398 15538 18450
rect 18734 18398 18786 18450
rect 20078 18398 20130 18450
rect 21310 18398 21362 18450
rect 22430 18398 22482 18450
rect 22654 18398 22706 18450
rect 23774 18398 23826 18450
rect 25454 18398 25506 18450
rect 27134 18398 27186 18450
rect 29150 18398 29202 18450
rect 29374 18398 29426 18450
rect 30382 18398 30434 18450
rect 35534 18398 35586 18450
rect 36542 18398 36594 18450
rect 37214 18398 37266 18450
rect 37774 18398 37826 18450
rect 38782 18398 38834 18450
rect 39230 18398 39282 18450
rect 39454 18398 39506 18450
rect 43262 18398 43314 18450
rect 43598 18398 43650 18450
rect 45838 18398 45890 18450
rect 49646 18398 49698 18450
rect 50542 18398 50594 18450
rect 6526 18286 6578 18338
rect 9774 18286 9826 18338
rect 14254 18286 14306 18338
rect 15262 18286 15314 18338
rect 17726 18286 17778 18338
rect 23326 18286 23378 18338
rect 25566 18286 25618 18338
rect 26014 18286 26066 18338
rect 27694 18286 27746 18338
rect 28030 18286 28082 18338
rect 35758 18286 35810 18338
rect 37438 18286 37490 18338
rect 38558 18286 38610 18338
rect 40126 18286 40178 18338
rect 46286 18286 46338 18338
rect 46846 18286 46898 18338
rect 47518 18286 47570 18338
rect 50318 18286 50370 18338
rect 5070 18174 5122 18226
rect 17390 18174 17442 18226
rect 23774 18174 23826 18226
rect 29934 18174 29986 18226
rect 31166 18174 31218 18226
rect 31502 18174 31554 18226
rect 36094 18174 36146 18226
rect 36990 18174 37042 18226
rect 38446 18174 38498 18226
rect 47406 18174 47458 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 9774 17838 9826 17890
rect 28254 17838 28306 17890
rect 34526 17838 34578 17890
rect 57934 17838 57986 17890
rect 4398 17726 4450 17778
rect 7758 17726 7810 17778
rect 8654 17726 8706 17778
rect 10670 17726 10722 17778
rect 11006 17726 11058 17778
rect 15822 17726 15874 17778
rect 23774 17726 23826 17778
rect 24782 17726 24834 17778
rect 31502 17726 31554 17778
rect 32622 17726 32674 17778
rect 34750 17726 34802 17778
rect 42142 17726 42194 17778
rect 45950 17726 46002 17778
rect 48750 17726 48802 17778
rect 5070 17614 5122 17666
rect 5742 17614 5794 17666
rect 7198 17614 7250 17666
rect 8318 17614 8370 17666
rect 10782 17614 10834 17666
rect 11342 17614 11394 17666
rect 13582 17614 13634 17666
rect 14590 17614 14642 17666
rect 15038 17614 15090 17666
rect 17614 17614 17666 17666
rect 17726 17614 17778 17666
rect 17950 17614 18002 17666
rect 18174 17614 18226 17666
rect 19070 17614 19122 17666
rect 19294 17614 19346 17666
rect 22094 17614 22146 17666
rect 23102 17614 23154 17666
rect 24334 17614 24386 17666
rect 25902 17614 25954 17666
rect 26910 17614 26962 17666
rect 27246 17614 27298 17666
rect 29486 17614 29538 17666
rect 29934 17614 29986 17666
rect 30382 17614 30434 17666
rect 31054 17614 31106 17666
rect 32174 17614 32226 17666
rect 32734 17614 32786 17666
rect 34302 17614 34354 17666
rect 36206 17614 36258 17666
rect 41694 17614 41746 17666
rect 42702 17614 42754 17666
rect 43934 17614 43986 17666
rect 45726 17614 45778 17666
rect 46510 17614 46562 17666
rect 47070 17614 47122 17666
rect 48078 17614 48130 17666
rect 48638 17614 48690 17666
rect 49198 17614 49250 17666
rect 49534 17614 49586 17666
rect 51326 17614 51378 17666
rect 55582 17614 55634 17666
rect 1710 17502 1762 17554
rect 6526 17502 6578 17554
rect 11230 17502 11282 17554
rect 12910 17502 12962 17554
rect 13918 17502 13970 17554
rect 16830 17502 16882 17554
rect 17054 17502 17106 17554
rect 18734 17502 18786 17554
rect 21422 17502 21474 17554
rect 21534 17502 21586 17554
rect 22542 17502 22594 17554
rect 29822 17502 29874 17554
rect 31726 17502 31778 17554
rect 33406 17502 33458 17554
rect 35758 17502 35810 17554
rect 43038 17502 43090 17554
rect 46846 17502 46898 17554
rect 50654 17502 50706 17554
rect 51102 17502 51154 17554
rect 51662 17502 51714 17554
rect 14478 17390 14530 17442
rect 20638 17390 20690 17442
rect 21198 17390 21250 17442
rect 23102 17390 23154 17442
rect 29710 17390 29762 17442
rect 38782 17390 38834 17442
rect 39118 17390 39170 17442
rect 43374 17390 43426 17442
rect 47406 17390 47458 17442
rect 51214 17390 51266 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 5182 17054 5234 17106
rect 5518 17054 5570 17106
rect 6078 17054 6130 17106
rect 6974 17054 7026 17106
rect 7758 17054 7810 17106
rect 8094 17054 8146 17106
rect 10110 17054 10162 17106
rect 10558 17054 10610 17106
rect 24782 17054 24834 17106
rect 25454 17054 25506 17106
rect 30942 17054 30994 17106
rect 41694 17054 41746 17106
rect 8654 16942 8706 16994
rect 16270 16942 16322 16994
rect 17726 16942 17778 16994
rect 17950 16942 18002 16994
rect 18622 16942 18674 16994
rect 20638 16942 20690 16994
rect 23774 16942 23826 16994
rect 27582 16942 27634 16994
rect 29262 16942 29314 16994
rect 32510 16942 32562 16994
rect 37662 16942 37714 16994
rect 41470 16942 41522 16994
rect 43822 16942 43874 16994
rect 50206 16942 50258 16994
rect 58158 16942 58210 16994
rect 7198 16830 7250 16882
rect 10782 16830 10834 16882
rect 11342 16830 11394 16882
rect 14366 16830 14418 16882
rect 15262 16830 15314 16882
rect 15486 16830 15538 16882
rect 16830 16830 16882 16882
rect 18510 16830 18562 16882
rect 18846 16830 18898 16882
rect 19518 16830 19570 16882
rect 20862 16830 20914 16882
rect 22766 16830 22818 16882
rect 24334 16830 24386 16882
rect 25790 16830 25842 16882
rect 26574 16830 26626 16882
rect 27134 16830 27186 16882
rect 27806 16830 27858 16882
rect 28702 16830 28754 16882
rect 30270 16830 30322 16882
rect 31838 16830 31890 16882
rect 33854 16830 33906 16882
rect 34078 16830 34130 16882
rect 34414 16830 34466 16882
rect 35422 16830 35474 16882
rect 36094 16830 36146 16882
rect 36430 16830 36482 16882
rect 36766 16830 36818 16882
rect 37550 16830 37602 16882
rect 41022 16830 41074 16882
rect 41806 16830 41858 16882
rect 41918 16830 41970 16882
rect 42478 16830 42530 16882
rect 43374 16830 43426 16882
rect 45726 16830 45778 16882
rect 46958 16830 47010 16882
rect 47182 16830 47234 16882
rect 51102 16830 51154 16882
rect 51774 16830 51826 16882
rect 53118 16830 53170 16882
rect 6190 16718 6242 16770
rect 6526 16718 6578 16770
rect 5182 16606 5234 16658
rect 11678 16718 11730 16770
rect 13470 16718 13522 16770
rect 14926 16718 14978 16770
rect 19406 16718 19458 16770
rect 25230 16718 25282 16770
rect 25454 16718 25506 16770
rect 35534 16718 35586 16770
rect 37886 16718 37938 16770
rect 42590 16718 42642 16770
rect 45950 16718 46002 16770
rect 50318 16718 50370 16770
rect 14814 16606 14866 16658
rect 19854 16606 19906 16658
rect 26798 16606 26850 16658
rect 35086 16606 35138 16658
rect 46846 16606 46898 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 4286 16270 4338 16322
rect 4958 16270 5010 16322
rect 10782 16270 10834 16322
rect 37886 16270 37938 16322
rect 41918 16270 41970 16322
rect 57934 16270 57986 16322
rect 4286 16158 4338 16210
rect 5182 16158 5234 16210
rect 9774 16158 9826 16210
rect 10334 16158 10386 16210
rect 15262 16158 15314 16210
rect 16494 16158 16546 16210
rect 17166 16158 17218 16210
rect 19742 16158 19794 16210
rect 23438 16158 23490 16210
rect 26910 16158 26962 16210
rect 29710 16158 29762 16210
rect 35982 16158 36034 16210
rect 51214 16158 51266 16210
rect 6974 16046 7026 16098
rect 7422 16046 7474 16098
rect 7534 16046 7586 16098
rect 7646 16046 7698 16098
rect 8878 16046 8930 16098
rect 10446 16046 10498 16098
rect 12350 16046 12402 16098
rect 13582 16046 13634 16098
rect 14478 16046 14530 16098
rect 15598 16046 15650 16098
rect 16830 16046 16882 16098
rect 17838 16046 17890 16098
rect 19966 16046 20018 16098
rect 20190 16046 20242 16098
rect 20526 16046 20578 16098
rect 21310 16046 21362 16098
rect 22430 16046 22482 16098
rect 23326 16046 23378 16098
rect 23998 16046 24050 16098
rect 25006 16046 25058 16098
rect 25902 16046 25954 16098
rect 26798 16046 26850 16098
rect 27806 16046 27858 16098
rect 29262 16046 29314 16098
rect 29822 16046 29874 16098
rect 33406 16046 33458 16098
rect 33518 16046 33570 16098
rect 34302 16046 34354 16098
rect 37438 16046 37490 16098
rect 38670 16046 38722 16098
rect 39902 16046 39954 16098
rect 40798 16046 40850 16098
rect 41246 16046 41298 16098
rect 41358 16046 41410 16098
rect 50206 16046 50258 16098
rect 50878 16046 50930 16098
rect 55582 16046 55634 16098
rect 4734 15934 4786 15986
rect 5854 15934 5906 15986
rect 13694 15934 13746 15986
rect 14590 15934 14642 15986
rect 15150 15934 15202 15986
rect 19854 15934 19906 15986
rect 20414 15934 20466 15986
rect 25118 15934 25170 15986
rect 25790 15934 25842 15986
rect 27022 15934 27074 15986
rect 27582 15934 27634 15986
rect 33630 15934 33682 15986
rect 34638 15934 34690 15986
rect 34862 15934 34914 15986
rect 35758 15934 35810 15986
rect 37102 15934 37154 15986
rect 38894 15934 38946 15986
rect 39230 15934 39282 15986
rect 39790 15934 39842 15986
rect 42030 15934 42082 15986
rect 42254 15934 42306 15986
rect 50094 15934 50146 15986
rect 51550 15934 51602 15986
rect 52670 15934 52722 15986
rect 53006 15934 53058 15986
rect 8094 15822 8146 15874
rect 14030 15822 14082 15874
rect 23886 15822 23938 15874
rect 29374 15822 29426 15874
rect 29598 15822 29650 15874
rect 30270 15822 30322 15874
rect 30830 15822 30882 15874
rect 31166 15822 31218 15874
rect 31614 15822 31666 15874
rect 33182 15822 33234 15874
rect 35198 15822 35250 15874
rect 38222 15822 38274 15874
rect 39006 15822 39058 15874
rect 42366 15822 42418 15874
rect 49870 15822 49922 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 5070 15486 5122 15538
rect 5518 15486 5570 15538
rect 5966 15486 6018 15538
rect 9550 15486 9602 15538
rect 10782 15486 10834 15538
rect 11230 15486 11282 15538
rect 17502 15486 17554 15538
rect 28142 15486 28194 15538
rect 29262 15486 29314 15538
rect 30158 15486 30210 15538
rect 40798 15486 40850 15538
rect 41022 15486 41074 15538
rect 43486 15486 43538 15538
rect 45054 15486 45106 15538
rect 45838 15486 45890 15538
rect 46846 15486 46898 15538
rect 7086 15374 7138 15426
rect 8430 15374 8482 15426
rect 11454 15374 11506 15426
rect 12014 15374 12066 15426
rect 19182 15374 19234 15426
rect 21422 15374 21474 15426
rect 22766 15374 22818 15426
rect 24670 15374 24722 15426
rect 26910 15374 26962 15426
rect 27694 15374 27746 15426
rect 31726 15374 31778 15426
rect 35310 15374 35362 15426
rect 45390 15374 45442 15426
rect 46734 15374 46786 15426
rect 47294 15374 47346 15426
rect 47630 15374 47682 15426
rect 48302 15374 48354 15426
rect 50990 15374 51042 15426
rect 51102 15374 51154 15426
rect 53342 15374 53394 15426
rect 7646 15262 7698 15314
rect 8990 15262 9042 15314
rect 11790 15262 11842 15314
rect 12574 15262 12626 15314
rect 14142 15262 14194 15314
rect 15486 15262 15538 15314
rect 18174 15262 18226 15314
rect 18734 15262 18786 15314
rect 20302 15262 20354 15314
rect 21870 15262 21922 15314
rect 22654 15262 22706 15314
rect 23774 15262 23826 15314
rect 25790 15262 25842 15314
rect 26574 15262 26626 15314
rect 28142 15262 28194 15314
rect 28702 15262 28754 15314
rect 28926 15262 28978 15314
rect 29598 15262 29650 15314
rect 31166 15262 31218 15314
rect 31614 15262 31666 15314
rect 32958 15262 33010 15314
rect 33406 15262 33458 15314
rect 33630 15262 33682 15314
rect 34414 15262 34466 15314
rect 34750 15262 34802 15314
rect 35086 15262 35138 15314
rect 37214 15262 37266 15314
rect 37438 15262 37490 15314
rect 37774 15262 37826 15314
rect 38110 15262 38162 15314
rect 38334 15262 38386 15314
rect 39006 15262 39058 15314
rect 39678 15262 39730 15314
rect 39790 15262 39842 15314
rect 41134 15262 41186 15314
rect 42142 15262 42194 15314
rect 42366 15262 42418 15314
rect 42478 15262 42530 15314
rect 43038 15262 43090 15314
rect 45614 15262 45666 15314
rect 46174 15262 46226 15314
rect 46510 15262 46562 15314
rect 47070 15262 47122 15314
rect 51326 15262 51378 15314
rect 51774 15262 51826 15314
rect 52670 15262 52722 15314
rect 53006 15262 53058 15314
rect 6414 15150 6466 15202
rect 9998 15150 10050 15202
rect 11902 15150 11954 15202
rect 13358 15150 13410 15202
rect 15598 15150 15650 15202
rect 18958 15150 19010 15202
rect 20190 15150 20242 15202
rect 22766 15150 22818 15202
rect 24222 15150 24274 15202
rect 25678 15150 25730 15202
rect 26350 15150 26402 15202
rect 29822 15150 29874 15202
rect 30718 15150 30770 15202
rect 33518 15150 33570 15202
rect 33966 15150 34018 15202
rect 34974 15150 35026 15202
rect 41582 15150 41634 15202
rect 45838 15150 45890 15202
rect 51886 15150 51938 15202
rect 15262 15038 15314 15090
rect 40238 15038 40290 15090
rect 42030 15038 42082 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 21870 14702 21922 14754
rect 33854 14702 33906 14754
rect 40126 14702 40178 14754
rect 49870 14702 49922 14754
rect 57934 14702 57986 14754
rect 5182 14590 5234 14642
rect 6638 14590 6690 14642
rect 7310 14590 7362 14642
rect 8318 14590 8370 14642
rect 12126 14590 12178 14642
rect 13582 14590 13634 14642
rect 20638 14590 20690 14642
rect 21982 14590 22034 14642
rect 28030 14590 28082 14642
rect 31502 14590 31554 14642
rect 36318 14590 36370 14642
rect 38558 14590 38610 14642
rect 39790 14590 39842 14642
rect 43822 14590 43874 14642
rect 45838 14590 45890 14642
rect 47070 14590 47122 14642
rect 6190 14478 6242 14530
rect 6974 14478 7026 14530
rect 7870 14478 7922 14530
rect 9662 14478 9714 14530
rect 11006 14478 11058 14530
rect 11678 14478 11730 14530
rect 12574 14478 12626 14530
rect 13694 14478 13746 14530
rect 15262 14478 15314 14530
rect 16606 14478 16658 14530
rect 17502 14478 17554 14530
rect 18174 14478 18226 14530
rect 20190 14478 20242 14530
rect 21534 14478 21586 14530
rect 22766 14478 22818 14530
rect 23550 14478 23602 14530
rect 23998 14478 24050 14530
rect 24334 14478 24386 14530
rect 25006 14478 25058 14530
rect 25230 14478 25282 14530
rect 26574 14478 26626 14530
rect 28478 14478 28530 14530
rect 31278 14478 31330 14530
rect 33182 14478 33234 14530
rect 34638 14478 34690 14530
rect 35086 14478 35138 14530
rect 35310 14478 35362 14530
rect 37886 14478 37938 14530
rect 38894 14478 38946 14530
rect 39454 14478 39506 14530
rect 41134 14478 41186 14530
rect 42142 14478 42194 14530
rect 42366 14478 42418 14530
rect 43150 14478 43202 14530
rect 44158 14478 44210 14530
rect 45390 14478 45442 14530
rect 48526 14478 48578 14530
rect 55582 14478 55634 14530
rect 8654 14366 8706 14418
rect 10894 14366 10946 14418
rect 11454 14366 11506 14418
rect 12014 14366 12066 14418
rect 13918 14366 13970 14418
rect 18734 14366 18786 14418
rect 22990 14366 23042 14418
rect 24782 14366 24834 14418
rect 26238 14366 26290 14418
rect 26910 14366 26962 14418
rect 27134 14366 27186 14418
rect 27806 14366 27858 14418
rect 30494 14366 30546 14418
rect 31726 14366 31778 14418
rect 33630 14366 33682 14418
rect 38670 14366 38722 14418
rect 41694 14366 41746 14418
rect 42254 14366 42306 14418
rect 42814 14366 42866 14418
rect 43262 14366 43314 14418
rect 45054 14366 45106 14418
rect 47518 14366 47570 14418
rect 17838 14254 17890 14306
rect 23326 14254 23378 14306
rect 23438 14254 23490 14306
rect 29486 14254 29538 14306
rect 35758 14254 35810 14306
rect 41470 14254 41522 14306
rect 41806 14254 41858 14306
rect 44830 14254 44882 14306
rect 44942 14254 44994 14306
rect 45726 14254 45778 14306
rect 45950 14254 46002 14306
rect 46174 14254 46226 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 6190 13918 6242 13970
rect 7422 13918 7474 13970
rect 7758 13918 7810 13970
rect 8878 13918 8930 13970
rect 9102 13918 9154 13970
rect 16942 13918 16994 13970
rect 21086 13918 21138 13970
rect 21310 13918 21362 13970
rect 25230 13918 25282 13970
rect 25902 13918 25954 13970
rect 31950 13918 32002 13970
rect 33294 13918 33346 13970
rect 44942 13918 44994 13970
rect 45166 13918 45218 13970
rect 47406 13918 47458 13970
rect 47630 13918 47682 13970
rect 51774 13918 51826 13970
rect 8318 13806 8370 13858
rect 8766 13806 8818 13858
rect 10558 13806 10610 13858
rect 20526 13806 20578 13858
rect 21534 13806 21586 13858
rect 23102 13806 23154 13858
rect 23998 13806 24050 13858
rect 24446 13806 24498 13858
rect 25566 13806 25618 13858
rect 27134 13806 27186 13858
rect 28142 13806 28194 13858
rect 30494 13806 30546 13858
rect 31054 13806 31106 13858
rect 33182 13806 33234 13858
rect 33630 13806 33682 13858
rect 35086 13806 35138 13858
rect 37774 13806 37826 13858
rect 38446 13806 38498 13858
rect 38670 13806 38722 13858
rect 39342 13806 39394 13858
rect 43486 13806 43538 13858
rect 43598 13806 43650 13858
rect 44830 13806 44882 13858
rect 45502 13806 45554 13858
rect 46734 13806 46786 13858
rect 52334 13806 52386 13858
rect 58158 13806 58210 13858
rect 6638 13694 6690 13746
rect 6862 13694 6914 13746
rect 7086 13694 7138 13746
rect 10222 13694 10274 13746
rect 11342 13694 11394 13746
rect 12686 13694 12738 13746
rect 13134 13694 13186 13746
rect 14926 13694 14978 13746
rect 15486 13694 15538 13746
rect 16270 13694 16322 13746
rect 17614 13694 17666 13746
rect 19182 13694 19234 13746
rect 20414 13694 20466 13746
rect 20974 13694 21026 13746
rect 21870 13694 21922 13746
rect 22990 13694 23042 13746
rect 23774 13694 23826 13746
rect 27022 13694 27074 13746
rect 28478 13694 28530 13746
rect 30270 13694 30322 13746
rect 30606 13694 30658 13746
rect 33854 13694 33906 13746
rect 34974 13694 35026 13746
rect 37326 13694 37378 13746
rect 39006 13694 39058 13746
rect 43262 13694 43314 13746
rect 45838 13694 45890 13746
rect 46398 13694 46450 13746
rect 47294 13694 47346 13746
rect 49870 13694 49922 13746
rect 50318 13694 50370 13746
rect 51326 13694 51378 13746
rect 51662 13694 51714 13746
rect 52222 13694 52274 13746
rect 10334 13582 10386 13634
rect 11006 13582 11058 13634
rect 18398 13582 18450 13634
rect 19406 13582 19458 13634
rect 22766 13582 22818 13634
rect 26014 13582 26066 13634
rect 28590 13582 28642 13634
rect 31390 13582 31442 13634
rect 34638 13582 34690 13634
rect 36990 13582 37042 13634
rect 45390 13582 45442 13634
rect 46846 13582 46898 13634
rect 50430 13582 50482 13634
rect 13246 13470 13298 13522
rect 16046 13470 16098 13522
rect 20078 13470 20130 13522
rect 31614 13470 31666 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 15150 13134 15202 13186
rect 17838 13134 17890 13186
rect 18958 13134 19010 13186
rect 25118 13134 25170 13186
rect 30830 13134 30882 13186
rect 31614 13134 31666 13186
rect 32510 13134 32562 13186
rect 42142 13134 42194 13186
rect 49534 13134 49586 13186
rect 50766 13134 50818 13186
rect 6526 13022 6578 13074
rect 7870 13022 7922 13074
rect 8654 13022 8706 13074
rect 10110 13022 10162 13074
rect 12126 13022 12178 13074
rect 12910 13022 12962 13074
rect 16606 13022 16658 13074
rect 17614 13022 17666 13074
rect 25230 13022 25282 13074
rect 27246 13022 27298 13074
rect 28702 13022 28754 13074
rect 32398 13022 32450 13074
rect 43486 13022 43538 13074
rect 48974 13022 49026 13074
rect 50206 13022 50258 13074
rect 6974 12910 7026 12962
rect 8094 12910 8146 12962
rect 8990 12910 9042 12962
rect 11342 12910 11394 12962
rect 11902 12910 11954 12962
rect 14030 12910 14082 12962
rect 16270 12910 16322 12962
rect 18846 12910 18898 12962
rect 19406 12910 19458 12962
rect 21758 12910 21810 12962
rect 22430 12910 22482 12962
rect 23550 12910 23602 12962
rect 24894 12910 24946 12962
rect 26462 12910 26514 12962
rect 26686 12910 26738 12962
rect 27582 12910 27634 12962
rect 28142 12910 28194 12962
rect 29374 12910 29426 12962
rect 32174 12910 32226 12962
rect 42030 12910 42082 12962
rect 42590 12910 42642 12962
rect 42814 12910 42866 12962
rect 49198 12910 49250 12962
rect 50094 12910 50146 12962
rect 7310 12798 7362 12850
rect 11230 12798 11282 12850
rect 12462 12798 12514 12850
rect 17390 12798 17442 12850
rect 19742 12798 19794 12850
rect 20190 12798 20242 12850
rect 29486 12798 29538 12850
rect 30046 12798 30098 12850
rect 36318 12798 36370 12850
rect 36430 12798 36482 12850
rect 41918 12798 41970 12850
rect 13694 12686 13746 12738
rect 20302 12686 20354 12738
rect 30382 12686 30434 12738
rect 31054 12686 31106 12738
rect 31502 12686 31554 12738
rect 35870 12686 35922 12738
rect 36094 12686 36146 12738
rect 41582 12686 41634 12738
rect 58158 12686 58210 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 8206 12350 8258 12402
rect 9998 12350 10050 12402
rect 13246 12350 13298 12402
rect 15486 12350 15538 12402
rect 16830 12350 16882 12402
rect 22542 12350 22594 12402
rect 22766 12350 22818 12402
rect 23102 12350 23154 12402
rect 24222 12350 24274 12402
rect 25454 12350 25506 12402
rect 26350 12350 26402 12402
rect 26686 12350 26738 12402
rect 27358 12350 27410 12402
rect 27806 12350 27858 12402
rect 28254 12350 28306 12402
rect 30830 12350 30882 12402
rect 33294 12350 33346 12402
rect 35198 12350 35250 12402
rect 38446 12350 38498 12402
rect 38782 12350 38834 12402
rect 50654 12350 50706 12402
rect 10222 12238 10274 12290
rect 11566 12238 11618 12290
rect 11790 12238 11842 12290
rect 14030 12238 14082 12290
rect 17950 12238 18002 12290
rect 21982 12238 22034 12290
rect 24446 12238 24498 12290
rect 26126 12238 26178 12290
rect 27694 12238 27746 12290
rect 29598 12238 29650 12290
rect 29710 12238 29762 12290
rect 30270 12238 30322 12290
rect 31054 12238 31106 12290
rect 31502 12238 31554 12290
rect 35870 12238 35922 12290
rect 47518 12238 47570 12290
rect 7310 12126 7362 12178
rect 7534 12126 7586 12178
rect 8766 12126 8818 12178
rect 11118 12126 11170 12178
rect 12350 12126 12402 12178
rect 13470 12126 13522 12178
rect 15262 12126 15314 12178
rect 18174 12126 18226 12178
rect 19630 12126 19682 12178
rect 21310 12126 21362 12178
rect 26014 12126 26066 12178
rect 29934 12126 29986 12178
rect 30494 12126 30546 12178
rect 33182 12126 33234 12178
rect 34750 12126 34802 12178
rect 35982 12126 36034 12178
rect 36878 12126 36930 12178
rect 39118 12126 39170 12178
rect 39678 12126 39730 12178
rect 42366 12126 42418 12178
rect 43374 12126 43426 12178
rect 44494 12126 44546 12178
rect 46622 12126 46674 12178
rect 50094 12126 50146 12178
rect 50318 12126 50370 12178
rect 6638 12014 6690 12066
rect 7086 12014 7138 12066
rect 10782 12014 10834 12066
rect 11902 12014 11954 12066
rect 17502 12014 17554 12066
rect 20414 12014 20466 12066
rect 23774 12014 23826 12066
rect 24334 12014 24386 12066
rect 28702 12014 28754 12066
rect 29262 12014 29314 12066
rect 33854 12014 33906 12066
rect 37214 12014 37266 12066
rect 41694 12014 41746 12066
rect 42590 12014 42642 12066
rect 43598 12014 43650 12066
rect 44046 12014 44098 12066
rect 46734 12014 46786 12066
rect 7870 11902 7922 11954
rect 10446 11902 10498 11954
rect 27806 11902 27858 11954
rect 31166 11902 31218 11954
rect 33294 11902 33346 11954
rect 36878 11902 36930 11954
rect 42030 11902 42082 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 22766 11566 22818 11618
rect 23550 11566 23602 11618
rect 24894 11566 24946 11618
rect 25454 11566 25506 11618
rect 46622 11566 46674 11618
rect 7534 11454 7586 11506
rect 15038 11454 15090 11506
rect 18398 11454 18450 11506
rect 20750 11454 20802 11506
rect 21758 11454 21810 11506
rect 24334 11454 24386 11506
rect 25678 11454 25730 11506
rect 31390 11454 31442 11506
rect 33742 11454 33794 11506
rect 37438 11454 37490 11506
rect 39678 11454 39730 11506
rect 41134 11454 41186 11506
rect 43822 11454 43874 11506
rect 45390 11454 45442 11506
rect 46398 11454 46450 11506
rect 46958 11454 47010 11506
rect 50206 11454 50258 11506
rect 57934 11454 57986 11506
rect 8430 11342 8482 11394
rect 9214 11342 9266 11394
rect 9774 11342 9826 11394
rect 10558 11342 10610 11394
rect 11902 11342 11954 11394
rect 12798 11342 12850 11394
rect 15262 11342 15314 11394
rect 16046 11342 16098 11394
rect 17054 11342 17106 11394
rect 17390 11342 17442 11394
rect 18958 11342 19010 11394
rect 19518 11342 19570 11394
rect 22094 11342 22146 11394
rect 22542 11342 22594 11394
rect 22990 11342 23042 11394
rect 23102 11342 23154 11394
rect 23774 11342 23826 11394
rect 23998 11342 24050 11394
rect 24222 11342 24274 11394
rect 25006 11342 25058 11394
rect 26462 11342 26514 11394
rect 27358 11342 27410 11394
rect 28590 11342 28642 11394
rect 29374 11342 29426 11394
rect 30158 11342 30210 11394
rect 31054 11342 31106 11394
rect 33294 11342 33346 11394
rect 34078 11342 34130 11394
rect 34750 11342 34802 11394
rect 35198 11342 35250 11394
rect 35310 11342 35362 11394
rect 36878 11342 36930 11394
rect 37326 11342 37378 11394
rect 37886 11342 37938 11394
rect 39454 11342 39506 11394
rect 40350 11342 40402 11394
rect 41806 11342 41858 11394
rect 42254 11342 42306 11394
rect 43374 11342 43426 11394
rect 43710 11342 43762 11394
rect 47294 11342 47346 11394
rect 47518 11342 47570 11394
rect 50318 11342 50370 11394
rect 55582 11342 55634 11394
rect 8878 11230 8930 11282
rect 12350 11230 12402 11282
rect 19854 11230 19906 11282
rect 19966 11230 20018 11282
rect 24446 11230 24498 11282
rect 26126 11230 26178 11282
rect 26462 11230 26514 11282
rect 27918 11230 27970 11282
rect 30270 11230 30322 11282
rect 30942 11230 30994 11282
rect 34526 11230 34578 11282
rect 37998 11230 38050 11282
rect 39790 11230 39842 11282
rect 42926 11230 42978 11282
rect 43934 11230 43986 11282
rect 50990 11230 51042 11282
rect 51326 11230 51378 11282
rect 51662 11230 51714 11282
rect 8094 11118 8146 11170
rect 11230 11118 11282 11170
rect 13806 11118 13858 11170
rect 20190 11118 20242 11170
rect 25790 11118 25842 11170
rect 26574 11118 26626 11170
rect 27582 11118 27634 11170
rect 32958 11118 33010 11170
rect 34974 11118 35026 11170
rect 37550 11118 37602 11170
rect 38222 11118 38274 11170
rect 41470 11118 41522 11170
rect 41694 11118 41746 11170
rect 42366 11118 42418 11170
rect 45838 11118 45890 11170
rect 47854 11118 47906 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 8206 10782 8258 10834
rect 8654 10782 8706 10834
rect 14254 10782 14306 10834
rect 16382 10782 16434 10834
rect 17614 10782 17666 10834
rect 17950 10782 18002 10834
rect 22990 10782 23042 10834
rect 23550 10782 23602 10834
rect 24110 10782 24162 10834
rect 24334 10782 24386 10834
rect 24446 10782 24498 10834
rect 28814 10782 28866 10834
rect 29262 10782 29314 10834
rect 30158 10782 30210 10834
rect 34750 10782 34802 10834
rect 36094 10782 36146 10834
rect 36318 10782 36370 10834
rect 9102 10670 9154 10722
rect 10222 10670 10274 10722
rect 14030 10670 14082 10722
rect 22542 10670 22594 10722
rect 25790 10670 25842 10722
rect 27134 10670 27186 10722
rect 31502 10670 31554 10722
rect 31838 10670 31890 10722
rect 33742 10670 33794 10722
rect 34190 10670 34242 10722
rect 34974 10670 35026 10722
rect 57710 10670 57762 10722
rect 10446 10558 10498 10610
rect 11454 10558 11506 10610
rect 12798 10558 12850 10610
rect 13470 10558 13522 10610
rect 15150 10558 15202 10610
rect 15374 10558 15426 10610
rect 15598 10558 15650 10610
rect 16830 10558 16882 10610
rect 18062 10558 18114 10610
rect 18958 10558 19010 10610
rect 19518 10558 19570 10610
rect 20750 10558 20802 10610
rect 21086 10558 21138 10610
rect 22206 10558 22258 10610
rect 23774 10558 23826 10610
rect 27022 10558 27074 10610
rect 28142 10558 28194 10610
rect 29934 10558 29986 10610
rect 30606 10558 30658 10610
rect 33518 10558 33570 10610
rect 35422 10558 35474 10610
rect 35982 10558 36034 10610
rect 37662 10558 37714 10610
rect 38558 10558 38610 10610
rect 39006 10558 39058 10610
rect 42142 10558 42194 10610
rect 42366 10558 42418 10610
rect 43038 10558 43090 10610
rect 46734 10558 46786 10610
rect 47630 10558 47682 10610
rect 48862 10558 48914 10610
rect 48974 10558 49026 10610
rect 10558 10446 10610 10498
rect 17950 10446 18002 10498
rect 19966 10446 20018 10498
rect 20302 10446 20354 10498
rect 21982 10446 22034 10498
rect 25342 10446 25394 10498
rect 26350 10446 26402 10498
rect 26910 10446 26962 10498
rect 30046 10446 30098 10498
rect 31278 10446 31330 10498
rect 34862 10446 34914 10498
rect 37886 10446 37938 10498
rect 39454 10446 39506 10498
rect 41246 10446 41298 10498
rect 41694 10446 41746 10498
rect 47070 10446 47122 10498
rect 58158 10446 58210 10498
rect 25230 10334 25282 10386
rect 26350 10334 26402 10386
rect 30942 10334 30994 10386
rect 33182 10334 33234 10386
rect 37326 10334 37378 10386
rect 41246 10334 41298 10386
rect 41694 10334 41746 10386
rect 50206 10334 50258 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 25454 9998 25506 10050
rect 25790 9998 25842 10050
rect 26462 9998 26514 10050
rect 34302 9998 34354 10050
rect 34638 9998 34690 10050
rect 48974 9998 49026 10050
rect 8542 9886 8594 9938
rect 9438 9886 9490 9938
rect 13582 9886 13634 9938
rect 14702 9886 14754 9938
rect 17054 9886 17106 9938
rect 19294 9886 19346 9938
rect 21758 9886 21810 9938
rect 23326 9886 23378 9938
rect 28478 9886 28530 9938
rect 29598 9886 29650 9938
rect 35870 9886 35922 9938
rect 40574 9886 40626 9938
rect 46286 9886 46338 9938
rect 47070 9886 47122 9938
rect 9774 9774 9826 9826
rect 10334 9774 10386 9826
rect 10894 9774 10946 9826
rect 11678 9774 11730 9826
rect 12238 9774 12290 9826
rect 13694 9774 13746 9826
rect 14926 9774 14978 9826
rect 15822 9774 15874 9826
rect 16830 9774 16882 9826
rect 17278 9774 17330 9826
rect 18174 9774 18226 9826
rect 19182 9774 19234 9826
rect 20190 9774 20242 9826
rect 20638 9774 20690 9826
rect 21310 9774 21362 9826
rect 21646 9774 21698 9826
rect 21870 9774 21922 9826
rect 22206 9774 22258 9826
rect 22766 9774 22818 9826
rect 23438 9774 23490 9826
rect 23774 9774 23826 9826
rect 24110 9774 24162 9826
rect 24446 9774 24498 9826
rect 26462 9774 26514 9826
rect 27022 9774 27074 9826
rect 27246 9774 27298 9826
rect 27470 9774 27522 9826
rect 27694 9774 27746 9826
rect 29150 9774 29202 9826
rect 33406 9774 33458 9826
rect 34078 9774 34130 9826
rect 38782 9774 38834 9826
rect 39118 9774 39170 9826
rect 39342 9774 39394 9826
rect 40014 9774 40066 9826
rect 40686 9774 40738 9826
rect 44046 9774 44098 9826
rect 44158 9774 44210 9826
rect 45054 9774 45106 9826
rect 46510 9774 46562 9826
rect 47182 9774 47234 9826
rect 8990 9662 9042 9714
rect 11566 9662 11618 9714
rect 14478 9662 14530 9714
rect 16718 9662 16770 9714
rect 18398 9662 18450 9714
rect 18846 9662 18898 9714
rect 19630 9662 19682 9714
rect 22542 9662 22594 9714
rect 24222 9662 24274 9714
rect 26126 9662 26178 9714
rect 34526 9662 34578 9714
rect 38446 9662 38498 9714
rect 38558 9662 38610 9714
rect 41358 9662 41410 9714
rect 45390 9662 45442 9714
rect 45838 9662 45890 9714
rect 47854 9662 47906 9714
rect 49198 9662 49250 9714
rect 9998 9550 10050 9602
rect 12126 9550 12178 9602
rect 13022 9550 13074 9602
rect 15486 9550 15538 9602
rect 19406 9550 19458 9602
rect 20526 9550 20578 9602
rect 20750 9550 20802 9602
rect 22654 9550 22706 9602
rect 23214 9550 23266 9602
rect 25118 9550 25170 9602
rect 25678 9550 25730 9602
rect 27358 9550 27410 9602
rect 32398 9550 32450 9602
rect 33518 9550 33570 9602
rect 33630 9550 33682 9602
rect 35758 9550 35810 9602
rect 38222 9550 38274 9602
rect 43822 9550 43874 9602
rect 44270 9550 44322 9602
rect 49086 9550 49138 9602
rect 58158 9550 58210 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 9998 9214 10050 9266
rect 10894 9214 10946 9266
rect 11790 9214 11842 9266
rect 14366 9214 14418 9266
rect 15822 9214 15874 9266
rect 16270 9214 16322 9266
rect 16382 9214 16434 9266
rect 18958 9214 19010 9266
rect 23214 9214 23266 9266
rect 24110 9214 24162 9266
rect 26014 9214 26066 9266
rect 26798 9214 26850 9266
rect 27134 9214 27186 9266
rect 27582 9214 27634 9266
rect 27918 9214 27970 9266
rect 28254 9214 28306 9266
rect 28814 9214 28866 9266
rect 36766 9214 36818 9266
rect 39790 9214 39842 9266
rect 40462 9214 40514 9266
rect 45390 9214 45442 9266
rect 51438 9214 51490 9266
rect 12126 9102 12178 9154
rect 13470 9102 13522 9154
rect 14926 9102 14978 9154
rect 18510 9102 18562 9154
rect 19406 9102 19458 9154
rect 24558 9102 24610 9154
rect 26574 9102 26626 9154
rect 29262 9102 29314 9154
rect 29710 9102 29762 9154
rect 36094 9102 36146 9154
rect 42590 9102 42642 9154
rect 49086 9102 49138 9154
rect 50542 9102 50594 9154
rect 50766 9102 50818 9154
rect 10446 8990 10498 9042
rect 12574 8990 12626 9042
rect 14814 8990 14866 9042
rect 15934 8990 15986 9042
rect 16494 8990 16546 9042
rect 16942 8990 16994 9042
rect 17950 8990 18002 9042
rect 18174 8990 18226 9042
rect 18734 8990 18786 9042
rect 19070 8990 19122 9042
rect 19294 8990 19346 9042
rect 21646 8990 21698 9042
rect 21982 8990 22034 9042
rect 22766 8990 22818 9042
rect 24446 8990 24498 9042
rect 24782 8990 24834 9042
rect 25566 8990 25618 9042
rect 25678 8990 25730 9042
rect 25902 8990 25954 9042
rect 26462 8990 26514 9042
rect 31614 8990 31666 9042
rect 31950 8990 32002 9042
rect 35310 8990 35362 9042
rect 35982 8990 36034 9042
rect 38670 8990 38722 9042
rect 39118 8990 39170 9042
rect 39342 8990 39394 9042
rect 39678 8990 39730 9042
rect 41806 8990 41858 9042
rect 42254 8990 42306 9042
rect 42814 8990 42866 9042
rect 43150 8990 43202 9042
rect 44494 8990 44546 9042
rect 44942 8990 44994 9042
rect 45614 8990 45666 9042
rect 45838 8990 45890 9042
rect 46174 8990 46226 9042
rect 49422 8990 49474 9042
rect 49982 8990 50034 9042
rect 11342 8878 11394 8930
rect 12686 8878 12738 8930
rect 13918 8878 13970 8930
rect 25790 8878 25842 8930
rect 32510 8878 32562 8930
rect 43038 8878 43090 8930
rect 46062 8878 46114 8930
rect 49198 8878 49250 8930
rect 51326 8878 51378 8930
rect 13358 8766 13410 8818
rect 17502 8766 17554 8818
rect 28814 8766 28866 8818
rect 29486 8766 29538 8818
rect 34974 8766 35026 8818
rect 39790 8766 39842 8818
rect 44718 8766 44770 8818
rect 50878 8766 50930 8818
rect 51214 8766 51266 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 14814 8430 14866 8482
rect 25006 8430 25058 8482
rect 45838 8430 45890 8482
rect 10894 8318 10946 8370
rect 11342 8318 11394 8370
rect 21422 8318 21474 8370
rect 27918 8318 27970 8370
rect 28254 8318 28306 8370
rect 35310 8318 35362 8370
rect 43150 8318 43202 8370
rect 45502 8318 45554 8370
rect 50542 8318 50594 8370
rect 57934 8318 57986 8370
rect 11566 8206 11618 8258
rect 13806 8206 13858 8258
rect 14366 8206 14418 8258
rect 14926 8206 14978 8258
rect 15262 8206 15314 8258
rect 15934 8206 15986 8258
rect 16270 8206 16322 8258
rect 16830 8206 16882 8258
rect 18510 8206 18562 8258
rect 20078 8206 20130 8258
rect 23326 8206 23378 8258
rect 23774 8206 23826 8258
rect 23998 8206 24050 8258
rect 24894 8206 24946 8258
rect 26910 8206 26962 8258
rect 29038 8206 29090 8258
rect 29486 8206 29538 8258
rect 32062 8206 32114 8258
rect 35534 8206 35586 8258
rect 41470 8206 41522 8258
rect 41918 8206 41970 8258
rect 42478 8206 42530 8258
rect 42590 8206 42642 8258
rect 45166 8206 45218 8258
rect 45390 8206 45442 8258
rect 48190 8206 48242 8258
rect 48526 8206 48578 8258
rect 49534 8206 49586 8258
rect 50878 8206 50930 8258
rect 55582 8206 55634 8258
rect 17502 8094 17554 8146
rect 18846 8094 18898 8146
rect 19966 8094 20018 8146
rect 27582 8094 27634 8146
rect 27806 8094 27858 8146
rect 28366 8094 28418 8146
rect 28478 8094 28530 8146
rect 29710 8094 29762 8146
rect 30046 8094 30098 8146
rect 30382 8094 30434 8146
rect 32174 8094 32226 8146
rect 32734 8094 32786 8146
rect 33070 8094 33122 8146
rect 36094 8094 36146 8146
rect 38670 8094 38722 8146
rect 42702 8094 42754 8146
rect 48638 8094 48690 8146
rect 51662 8094 51714 8146
rect 51998 8094 52050 8146
rect 11902 7982 11954 8034
rect 12238 7982 12290 8034
rect 12574 7982 12626 8034
rect 16046 7982 16098 8034
rect 25902 7982 25954 8034
rect 26350 7982 26402 8034
rect 27246 7982 27298 8034
rect 29598 7982 29650 8034
rect 30158 7982 30210 8034
rect 33182 7982 33234 8034
rect 33406 7982 33458 8034
rect 38782 7982 38834 8034
rect 39006 7982 39058 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 9886 7646 9938 7698
rect 15374 7646 15426 7698
rect 16942 7646 16994 7698
rect 17838 7646 17890 7698
rect 19854 7646 19906 7698
rect 20078 7646 20130 7698
rect 21534 7646 21586 7698
rect 21870 7646 21922 7698
rect 22542 7646 22594 7698
rect 22990 7646 23042 7698
rect 23438 7646 23490 7698
rect 23886 7646 23938 7698
rect 27358 7646 27410 7698
rect 27806 7646 27858 7698
rect 28254 7646 28306 7698
rect 35534 7646 35586 7698
rect 36094 7646 36146 7698
rect 58158 7646 58210 7698
rect 12238 7534 12290 7586
rect 14590 7534 14642 7586
rect 16382 7534 16434 7586
rect 17614 7534 17666 7586
rect 20190 7534 20242 7586
rect 25342 7534 25394 7586
rect 26014 7534 26066 7586
rect 32510 7534 32562 7586
rect 33406 7534 33458 7586
rect 34414 7534 34466 7586
rect 48974 7534 49026 7586
rect 51326 7534 51378 7586
rect 10222 7422 10274 7474
rect 10670 7422 10722 7474
rect 11006 7422 11058 7474
rect 12014 7422 12066 7474
rect 13470 7422 13522 7474
rect 15486 7422 15538 7474
rect 15934 7422 15986 7474
rect 16046 7422 16098 7474
rect 18622 7422 18674 7474
rect 19294 7422 19346 7474
rect 20638 7422 20690 7474
rect 20862 7422 20914 7474
rect 21646 7422 21698 7474
rect 21982 7422 22034 7474
rect 24222 7422 24274 7474
rect 24558 7422 24610 7474
rect 25678 7422 25730 7474
rect 26238 7422 26290 7474
rect 28926 7422 28978 7474
rect 30046 7422 30098 7474
rect 32062 7422 32114 7474
rect 33966 7422 34018 7474
rect 34862 7422 34914 7474
rect 35310 7422 35362 7474
rect 35646 7422 35698 7474
rect 42254 7422 42306 7474
rect 42814 7422 42866 7474
rect 43374 7422 43426 7474
rect 43934 7422 43986 7474
rect 45502 7422 45554 7474
rect 45838 7422 45890 7474
rect 49310 7422 49362 7474
rect 50878 7422 50930 7474
rect 51214 7422 51266 7474
rect 16270 7310 16322 7362
rect 17950 7310 18002 7362
rect 18510 7310 18562 7362
rect 19406 7310 19458 7362
rect 24670 7310 24722 7362
rect 26014 7310 26066 7362
rect 28814 7310 28866 7362
rect 31950 7310 32002 7362
rect 34638 7310 34690 7362
rect 42142 7310 42194 7362
rect 47070 7310 47122 7362
rect 49422 7310 49474 7362
rect 21086 7198 21138 7250
rect 22430 7198 22482 7250
rect 23102 7198 23154 7250
rect 24334 7198 24386 7250
rect 29822 7198 29874 7250
rect 43598 7198 43650 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 14030 6862 14082 6914
rect 14702 6862 14754 6914
rect 18174 6862 18226 6914
rect 25006 6862 25058 6914
rect 35870 6862 35922 6914
rect 39118 6862 39170 6914
rect 9886 6750 9938 6802
rect 14478 6750 14530 6802
rect 16158 6750 16210 6802
rect 19966 6750 20018 6802
rect 23102 6750 23154 6802
rect 24894 6750 24946 6802
rect 28366 6750 28418 6802
rect 29262 6750 29314 6802
rect 38558 6750 38610 6802
rect 48302 6750 48354 6802
rect 11678 6638 11730 6690
rect 12238 6638 12290 6690
rect 12798 6638 12850 6690
rect 13806 6638 13858 6690
rect 14254 6638 14306 6690
rect 15038 6638 15090 6690
rect 15822 6638 15874 6690
rect 16606 6638 16658 6690
rect 18398 6638 18450 6690
rect 19294 6638 19346 6690
rect 19630 6638 19682 6690
rect 20190 6638 20242 6690
rect 21422 6638 21474 6690
rect 22654 6638 22706 6690
rect 23998 6638 24050 6690
rect 24670 6638 24722 6690
rect 25342 6638 25394 6690
rect 26798 6638 26850 6690
rect 27470 6638 27522 6690
rect 28478 6638 28530 6690
rect 31390 6638 31442 6690
rect 31614 6638 31666 6690
rect 32062 6638 32114 6690
rect 32622 6638 32674 6690
rect 33966 6638 34018 6690
rect 35198 6638 35250 6690
rect 36990 6638 37042 6690
rect 38110 6638 38162 6690
rect 38670 6638 38722 6690
rect 39006 6638 39058 6690
rect 47854 6638 47906 6690
rect 49086 6638 49138 6690
rect 11342 6526 11394 6578
rect 19854 6526 19906 6578
rect 20414 6526 20466 6578
rect 20750 6526 20802 6578
rect 24446 6526 24498 6578
rect 26350 6526 26402 6578
rect 28142 6526 28194 6578
rect 35086 6526 35138 6578
rect 11902 6414 11954 6466
rect 15150 6414 15202 6466
rect 15486 6414 15538 6466
rect 15710 6414 15762 6466
rect 20638 6414 20690 6466
rect 22094 6414 22146 6466
rect 22318 6414 22370 6466
rect 25566 6414 25618 6466
rect 26462 6414 26514 6466
rect 31502 6414 31554 6466
rect 37326 6414 37378 6466
rect 38446 6414 38498 6466
rect 39118 6414 39170 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 12350 6078 12402 6130
rect 12686 6078 12738 6130
rect 13694 6078 13746 6130
rect 14254 6078 14306 6130
rect 18622 6078 18674 6130
rect 18958 6078 19010 6130
rect 20190 6078 20242 6130
rect 21534 6078 21586 6130
rect 22094 6078 22146 6130
rect 23326 6078 23378 6130
rect 23662 6078 23714 6130
rect 25342 6078 25394 6130
rect 25454 6078 25506 6130
rect 26686 6078 26738 6130
rect 26910 6078 26962 6130
rect 29934 6078 29986 6130
rect 30606 6078 30658 6130
rect 39902 6078 39954 6130
rect 41358 6078 41410 6130
rect 42254 6078 42306 6130
rect 44270 6078 44322 6130
rect 15262 5966 15314 6018
rect 17726 5966 17778 6018
rect 19854 5966 19906 6018
rect 20638 5966 20690 6018
rect 22654 5966 22706 6018
rect 24334 5966 24386 6018
rect 24782 5966 24834 6018
rect 28030 5966 28082 6018
rect 29822 5966 29874 6018
rect 31502 5966 31554 6018
rect 31614 5966 31666 6018
rect 35870 5966 35922 6018
rect 37438 5966 37490 6018
rect 48750 5966 48802 6018
rect 48862 5966 48914 6018
rect 50990 5966 51042 6018
rect 15486 5854 15538 5906
rect 16270 5854 16322 5906
rect 17838 5854 17890 5906
rect 18286 5854 18338 5906
rect 18510 5854 18562 5906
rect 19518 5854 19570 5906
rect 20526 5854 20578 5906
rect 21646 5854 21698 5906
rect 22990 5854 23042 5906
rect 25230 5854 25282 5906
rect 25902 5854 25954 5906
rect 26350 5854 26402 5906
rect 27134 5854 27186 5906
rect 28142 5854 28194 5906
rect 29038 5854 29090 5906
rect 31838 5854 31890 5906
rect 36206 5854 36258 5906
rect 38446 5854 38498 5906
rect 39118 5854 39170 5906
rect 39678 5854 39730 5906
rect 40798 5854 40850 5906
rect 41246 5854 41298 5906
rect 41470 5854 41522 5906
rect 41694 5854 41746 5906
rect 42142 5854 42194 5906
rect 42366 5854 42418 5906
rect 43150 5854 43202 5906
rect 43486 5854 43538 5906
rect 44158 5854 44210 5906
rect 44606 5854 44658 5906
rect 46734 5854 46786 5906
rect 47630 5854 47682 5906
rect 49422 5854 49474 5906
rect 49646 5854 49698 5906
rect 50318 5854 50370 5906
rect 50654 5854 50706 5906
rect 11902 5742 11954 5794
rect 13134 5742 13186 5794
rect 13806 5742 13858 5794
rect 14814 5742 14866 5794
rect 16158 5742 16210 5794
rect 22766 5742 22818 5794
rect 27022 5742 27074 5794
rect 27806 5742 27858 5794
rect 29374 5742 29426 5794
rect 37662 5742 37714 5794
rect 40014 5742 40066 5794
rect 43262 5742 43314 5794
rect 45166 5742 45218 5794
rect 46398 5742 46450 5794
rect 47294 5742 47346 5794
rect 13470 5630 13522 5682
rect 14590 5630 14642 5682
rect 16494 5630 16546 5682
rect 29934 5630 29986 5682
rect 38334 5630 38386 5682
rect 42926 5630 42978 5682
rect 43710 5630 43762 5682
rect 44382 5630 44434 5682
rect 45278 5630 45330 5682
rect 47854 5630 47906 5682
rect 48190 5630 48242 5682
rect 48862 5630 48914 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 14814 5294 14866 5346
rect 15486 5294 15538 5346
rect 19854 5294 19906 5346
rect 20526 5294 20578 5346
rect 34750 5294 34802 5346
rect 39678 5294 39730 5346
rect 39902 5294 39954 5346
rect 40574 5294 40626 5346
rect 40798 5294 40850 5346
rect 44158 5294 44210 5346
rect 13022 5182 13074 5234
rect 13694 5182 13746 5234
rect 14030 5182 14082 5234
rect 14590 5182 14642 5234
rect 16270 5182 16322 5234
rect 22430 5182 22482 5234
rect 23886 5182 23938 5234
rect 24334 5182 24386 5234
rect 25118 5182 25170 5234
rect 25678 5182 25730 5234
rect 26910 5182 26962 5234
rect 41582 5238 41634 5290
rect 46398 5294 46450 5346
rect 27694 5182 27746 5234
rect 28142 5182 28194 5234
rect 30382 5182 30434 5234
rect 32734 5182 32786 5234
rect 40350 5182 40402 5234
rect 43262 5182 43314 5234
rect 46734 5182 46786 5234
rect 48078 5182 48130 5234
rect 15150 5070 15202 5122
rect 15486 5070 15538 5122
rect 16942 5070 16994 5122
rect 17614 5070 17666 5122
rect 17838 5070 17890 5122
rect 17950 5070 18002 5122
rect 18398 5070 18450 5122
rect 18622 5070 18674 5122
rect 18958 5070 19010 5122
rect 19742 5070 19794 5122
rect 21758 5070 21810 5122
rect 21982 5070 22034 5122
rect 22206 5070 22258 5122
rect 22654 5070 22706 5122
rect 24782 5070 24834 5122
rect 25454 5070 25506 5122
rect 25902 5070 25954 5122
rect 26014 5070 26066 5122
rect 26350 5070 26402 5122
rect 27022 5070 27074 5122
rect 28478 5070 28530 5122
rect 29150 5070 29202 5122
rect 32174 5070 32226 5122
rect 32846 5070 32898 5122
rect 33966 5070 34018 5122
rect 34526 5070 34578 5122
rect 38446 5070 38498 5122
rect 38670 5070 38722 5122
rect 39454 5070 39506 5122
rect 41246 5070 41298 5122
rect 41806 5070 41858 5122
rect 43038 5070 43090 5122
rect 45390 5070 45442 5122
rect 45950 5070 46002 5122
rect 46062 5070 46114 5122
rect 47070 5070 47122 5122
rect 48526 5070 48578 5122
rect 49086 5070 49138 5122
rect 49534 5070 49586 5122
rect 50094 5070 50146 5122
rect 15822 4958 15874 5010
rect 16606 4958 16658 5010
rect 19182 4958 19234 5010
rect 19518 4958 19570 5010
rect 20750 4958 20802 5010
rect 21422 4958 21474 5010
rect 26798 4958 26850 5010
rect 29374 4958 29426 5010
rect 29710 4958 29762 5010
rect 31838 4958 31890 5010
rect 33182 4958 33234 5010
rect 34078 4958 34130 5010
rect 34302 4958 34354 5010
rect 35646 4958 35698 5010
rect 38894 4958 38946 5010
rect 40014 4958 40066 5010
rect 42142 4958 42194 5010
rect 43710 4958 43762 5010
rect 44046 4958 44098 5010
rect 46510 4958 46562 5010
rect 48414 4958 48466 5010
rect 50430 4958 50482 5010
rect 51214 4958 51266 5010
rect 51326 4958 51378 5010
rect 14926 4846 14978 4898
rect 19070 4846 19122 4898
rect 20190 4846 20242 4898
rect 21534 4846 21586 4898
rect 22766 4846 22818 4898
rect 22878 4846 22930 4898
rect 35086 4846 35138 4898
rect 35310 4846 35362 4898
rect 35534 4846 35586 4898
rect 44158 4846 44210 4898
rect 47406 4846 47458 4898
rect 49422 4846 49474 4898
rect 49646 4846 49698 4898
rect 50766 4846 50818 4898
rect 50990 4846 51042 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 14366 4510 14418 4562
rect 15262 4510 15314 4562
rect 15598 4510 15650 4562
rect 16942 4510 16994 4562
rect 17614 4510 17666 4562
rect 18398 4510 18450 4562
rect 19966 4510 20018 4562
rect 21086 4510 21138 4562
rect 21870 4510 21922 4562
rect 23774 4510 23826 4562
rect 24334 4510 24386 4562
rect 24670 4510 24722 4562
rect 25454 4510 25506 4562
rect 26238 4510 26290 4562
rect 27246 4510 27298 4562
rect 28814 4510 28866 4562
rect 29486 4510 29538 4562
rect 30382 4510 30434 4562
rect 30718 4510 30770 4562
rect 30830 4510 30882 4562
rect 33070 4510 33122 4562
rect 34078 4510 34130 4562
rect 39566 4510 39618 4562
rect 42926 4510 42978 4562
rect 46846 4510 46898 4562
rect 50654 4510 50706 4562
rect 18846 4398 18898 4450
rect 19070 4398 19122 4450
rect 19294 4398 19346 4450
rect 22206 4398 22258 4450
rect 22430 4398 22482 4450
rect 23438 4398 23490 4450
rect 25230 4398 25282 4450
rect 28926 4398 28978 4450
rect 32286 4398 32338 4450
rect 33630 4398 33682 4450
rect 34526 4398 34578 4450
rect 39006 4398 39058 4450
rect 39342 4398 39394 4450
rect 42814 4398 42866 4450
rect 43598 4398 43650 4450
rect 49086 4398 49138 4450
rect 50766 4398 50818 4450
rect 19854 4286 19906 4338
rect 22766 4286 22818 4338
rect 30606 4286 30658 4338
rect 31838 4286 31890 4338
rect 33406 4286 33458 4338
rect 34302 4286 34354 4338
rect 35086 4286 35138 4338
rect 38558 4286 38610 4338
rect 43374 4286 43426 4338
rect 43934 4286 43986 4338
rect 47406 4286 47458 4338
rect 51326 4286 51378 4338
rect 14702 4174 14754 4226
rect 16494 4174 16546 4226
rect 19630 4174 19682 4226
rect 20526 4174 20578 4226
rect 21534 4174 21586 4226
rect 25566 4174 25618 4226
rect 31390 4174 31442 4226
rect 34414 4174 34466 4226
rect 35310 4174 35362 4226
rect 38110 4174 38162 4226
rect 39678 4174 39730 4226
rect 48862 4174 48914 4226
rect 16494 4062 16546 4114
rect 16718 4062 16770 4114
rect 22318 4062 22370 4114
rect 22990 4062 23042 4114
rect 28814 4062 28866 4114
rect 35870 4062 35922 4114
rect 44942 4062 44994 4114
rect 47182 4062 47234 4114
rect 52334 4062 52386 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 17054 3726 17106 3778
rect 18174 3726 18226 3778
rect 20750 3726 20802 3778
rect 21310 3726 21362 3778
rect 14926 3614 14978 3666
rect 15374 3614 15426 3666
rect 15822 3614 15874 3666
rect 16494 3614 16546 3666
rect 17278 3614 17330 3666
rect 17726 3614 17778 3666
rect 18174 3614 18226 3666
rect 18622 3614 18674 3666
rect 19742 3614 19794 3666
rect 20190 3614 20242 3666
rect 20974 3614 21026 3666
rect 21310 3614 21362 3666
rect 22990 3614 23042 3666
rect 23438 3614 23490 3666
rect 28814 3614 28866 3666
rect 32958 3614 33010 3666
rect 44606 3614 44658 3666
rect 52222 3614 52274 3666
rect 19294 3502 19346 3554
rect 21982 3502 22034 3554
rect 29038 3502 29090 3554
rect 32174 3502 32226 3554
rect 33070 3502 33122 3554
rect 38558 3502 38610 3554
rect 38894 3502 38946 3554
rect 44046 3502 44098 3554
rect 47518 3502 47570 3554
rect 51438 3502 51490 3554
rect 38670 3390 38722 3442
rect 48974 3390 49026 3442
rect 5518 3278 5570 3330
rect 9662 3278 9714 3330
rect 30046 3278 30098 3330
rect 54126 3278 54178 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
<< metal2 >>
rect 5376 59200 5488 60000
rect 6048 59200 6160 60000
rect 7392 59200 7504 60000
rect 8736 59200 8848 60000
rect 9408 59200 9520 60000
rect 10752 59200 10864 60000
rect 11424 59200 11536 60000
rect 30912 59200 31024 60000
rect 40992 59200 41104 60000
rect 45696 59200 45808 60000
rect 52416 59200 52528 60000
rect 54432 59200 54544 60000
rect 55104 59200 55216 60000
rect 5404 56308 5460 59200
rect 5628 56308 5684 56318
rect 5404 56306 5684 56308
rect 5404 56254 5630 56306
rect 5682 56254 5684 56306
rect 5404 56252 5684 56254
rect 6076 56308 6132 59200
rect 6300 56308 6356 56318
rect 6076 56306 6356 56308
rect 6076 56254 6302 56306
rect 6354 56254 6356 56306
rect 6076 56252 6356 56254
rect 7420 56308 7476 59200
rect 7644 56308 7700 56318
rect 7420 56306 7700 56308
rect 7420 56254 7646 56306
rect 7698 56254 7700 56306
rect 7420 56252 7700 56254
rect 5628 56242 5684 56252
rect 6300 56242 6356 56252
rect 7644 56242 7700 56252
rect 8764 55970 8820 59200
rect 9436 56308 9492 59200
rect 9660 56308 9716 56318
rect 9436 56306 9716 56308
rect 9436 56254 9662 56306
rect 9714 56254 9716 56306
rect 9436 56252 9716 56254
rect 10780 56308 10836 59200
rect 11004 56308 11060 56318
rect 10780 56306 11060 56308
rect 10780 56254 11006 56306
rect 11058 56254 11060 56306
rect 10780 56252 11060 56254
rect 11452 56308 11508 59200
rect 26684 57876 26740 57886
rect 15036 57764 15092 57774
rect 11676 56308 11732 56318
rect 11452 56306 11732 56308
rect 11452 56254 11678 56306
rect 11730 56254 11732 56306
rect 11452 56252 11732 56254
rect 9660 56242 9716 56252
rect 11004 56242 11060 56252
rect 11676 56242 11732 56252
rect 13804 56196 13860 56206
rect 13804 56102 13860 56140
rect 8764 55918 8766 55970
rect 8818 55918 8820 55970
rect 8764 55906 8820 55918
rect 12572 56084 12628 56094
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 1932 55410 1988 55422
rect 1932 55358 1934 55410
rect 1986 55358 1988 55410
rect 1932 54516 1988 55358
rect 4172 55298 4228 55310
rect 4172 55246 4174 55298
rect 4226 55246 4228 55298
rect 4172 55076 4228 55246
rect 4172 55010 4228 55020
rect 4732 55076 4788 55086
rect 4732 54982 4788 55020
rect 12460 55076 12516 55086
rect 1932 54450 1988 54460
rect 12012 54740 12068 54750
rect 11340 54404 11396 54414
rect 11900 54404 11956 54414
rect 11340 54402 11508 54404
rect 11340 54350 11342 54402
rect 11394 54350 11508 54402
rect 11340 54348 11508 54350
rect 11340 54338 11396 54348
rect 6524 54180 6580 54190
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 1708 51490 1764 51502
rect 1708 51438 1710 51490
rect 1762 51438 1764 51490
rect 1708 51156 1764 51438
rect 1708 51090 1764 51100
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 6524 50428 6580 54124
rect 9548 53730 9604 53742
rect 9548 53678 9550 53730
rect 9602 53678 9604 53730
rect 8316 53508 8372 53518
rect 8092 52276 8148 52286
rect 8316 52276 8372 53452
rect 8764 52276 8820 52286
rect 8092 52274 8372 52276
rect 8092 52222 8094 52274
rect 8146 52222 8372 52274
rect 8092 52220 8372 52222
rect 8092 52210 8148 52220
rect 8316 52162 8372 52220
rect 8652 52220 8764 52276
rect 8316 52110 8318 52162
rect 8370 52110 8372 52162
rect 8316 52098 8372 52110
rect 8540 52164 8596 52174
rect 6412 50372 6580 50428
rect 8204 51380 8260 51390
rect 8204 50482 8260 51324
rect 8204 50430 8206 50482
rect 8258 50430 8260 50482
rect 8204 50418 8260 50430
rect 7868 50372 7924 50382
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 1932 49138 1988 49150
rect 1932 49086 1934 49138
rect 1986 49086 1988 49138
rect 1932 48468 1988 49086
rect 4284 49026 4340 49038
rect 4284 48974 4286 49026
rect 4338 48974 4340 49026
rect 4284 48804 4340 48974
rect 4284 48738 4340 48748
rect 4732 48804 4788 48814
rect 4732 48710 4788 48748
rect 5628 48804 5684 48814
rect 1932 48402 1988 48412
rect 4284 48242 4340 48254
rect 4284 48190 4286 48242
rect 4338 48190 4340 48242
rect 1932 48020 1988 48030
rect 1932 47926 1988 47964
rect 4284 47348 4340 48190
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 4284 47282 4340 47292
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 1708 42866 1764 42878
rect 1708 42814 1710 42866
rect 1762 42814 1764 42866
rect 1708 42420 1764 42814
rect 1708 42354 1764 42364
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 1708 41300 1764 41310
rect 1708 41206 1764 41244
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 1708 39394 1764 39406
rect 1708 39342 1710 39394
rect 1762 39342 1764 39394
rect 1708 39060 1764 39342
rect 1708 38994 1764 39004
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 1708 37378 1764 37390
rect 1708 37326 1710 37378
rect 1762 37326 1764 37378
rect 1708 35700 1764 37326
rect 4284 37268 4340 37278
rect 2156 37044 2212 37054
rect 2156 36950 2212 36988
rect 1932 36596 1988 36606
rect 1932 36502 1988 36540
rect 4284 36482 4340 37212
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4284 36430 4286 36482
rect 4338 36430 4340 36482
rect 4284 36418 4340 36430
rect 1708 35634 1764 35644
rect 4284 35700 4340 35710
rect 4284 35606 4340 35644
rect 5516 35588 5572 35598
rect 1932 35474 1988 35486
rect 1932 35422 1934 35474
rect 1986 35422 1988 35474
rect 1932 35028 1988 35422
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 5516 35138 5572 35532
rect 5516 35086 5518 35138
rect 5570 35086 5572 35138
rect 5516 35074 5572 35086
rect 1932 34962 1988 34972
rect 5628 34468 5684 48748
rect 6076 45890 6132 45902
rect 6076 45838 6078 45890
rect 6130 45838 6132 45890
rect 6076 45668 6132 45838
rect 6300 45780 6356 45790
rect 6300 45686 6356 45724
rect 6076 45602 6132 45612
rect 6412 36932 6468 50372
rect 7420 50370 7924 50372
rect 7420 50318 7870 50370
rect 7922 50318 7924 50370
rect 7420 50316 7924 50318
rect 7420 49026 7476 50316
rect 7868 50306 7924 50316
rect 8540 50034 8596 52108
rect 8540 49982 8542 50034
rect 8594 49982 8596 50034
rect 8540 49970 8596 49982
rect 8316 49812 8372 49822
rect 8316 49718 8372 49756
rect 7420 48974 7422 49026
rect 7474 48974 7476 49026
rect 7420 47682 7476 48974
rect 7868 49026 7924 49038
rect 7868 48974 7870 49026
rect 7922 48974 7924 49026
rect 7868 48804 7924 48974
rect 7868 48738 7924 48748
rect 8204 48914 8260 48926
rect 8204 48862 8206 48914
rect 8258 48862 8260 48914
rect 8092 48468 8148 48478
rect 8092 48374 8148 48412
rect 7980 48244 8036 48254
rect 8204 48244 8260 48862
rect 7980 48242 8260 48244
rect 7980 48190 7982 48242
rect 8034 48190 8260 48242
rect 7980 48188 8260 48190
rect 7644 48132 7700 48142
rect 7644 48130 7812 48132
rect 7644 48078 7646 48130
rect 7698 48078 7812 48130
rect 7644 48076 7812 48078
rect 7644 48066 7700 48076
rect 7420 47630 7422 47682
rect 7474 47630 7476 47682
rect 7420 47618 7476 47630
rect 7308 47348 7364 47358
rect 7308 47068 7364 47292
rect 7084 47012 7364 47068
rect 6748 46786 6804 46798
rect 6748 46734 6750 46786
rect 6802 46734 6804 46786
rect 6524 45668 6580 45678
rect 6636 45668 6692 45678
rect 6748 45668 6804 46734
rect 7084 46674 7140 47012
rect 7084 46622 7086 46674
rect 7138 46622 7140 46674
rect 6972 46564 7028 46574
rect 7084 46564 7140 46622
rect 7028 46508 7140 46564
rect 6972 46498 7028 46508
rect 7644 46452 7700 46462
rect 7196 45892 7252 45902
rect 7196 45798 7252 45836
rect 7644 45890 7700 46396
rect 7644 45838 7646 45890
rect 7698 45838 7700 45890
rect 6580 45666 6804 45668
rect 6580 45614 6638 45666
rect 6690 45614 6804 45666
rect 6580 45612 6804 45614
rect 7644 45780 7700 45838
rect 6524 41188 6580 45612
rect 6636 45602 6692 45612
rect 7308 45106 7364 45118
rect 7308 45054 7310 45106
rect 7362 45054 7364 45106
rect 7308 44210 7364 45054
rect 7532 44548 7588 44558
rect 7644 44548 7700 45724
rect 7756 44996 7812 48076
rect 7868 44996 7924 45006
rect 7756 44940 7868 44996
rect 7868 44902 7924 44940
rect 7532 44546 7700 44548
rect 7532 44494 7534 44546
rect 7586 44494 7700 44546
rect 7532 44492 7700 44494
rect 7532 44482 7588 44492
rect 7308 44158 7310 44210
rect 7362 44158 7364 44210
rect 6972 43764 7028 43774
rect 7308 43764 7364 44158
rect 6972 43762 7588 43764
rect 6972 43710 6974 43762
rect 7026 43710 7588 43762
rect 6972 43708 7588 43710
rect 6972 43698 7028 43708
rect 6636 43540 6692 43550
rect 6636 43446 6692 43484
rect 7420 43538 7476 43550
rect 7420 43486 7422 43538
rect 7474 43486 7476 43538
rect 7308 42754 7364 42766
rect 7308 42702 7310 42754
rect 7362 42702 7364 42754
rect 7308 41748 7364 42702
rect 6636 41188 6692 41198
rect 6524 41132 6636 41188
rect 6636 41122 6692 41132
rect 7084 41188 7140 41198
rect 6860 40852 6916 40862
rect 6636 39620 6692 39630
rect 6636 39526 6692 39564
rect 6860 39506 6916 40796
rect 7084 40628 7140 41132
rect 7308 41074 7364 41692
rect 7308 41022 7310 41074
rect 7362 41022 7364 41074
rect 7196 40628 7252 40638
rect 7084 40626 7252 40628
rect 7084 40574 7198 40626
rect 7250 40574 7252 40626
rect 7084 40572 7252 40574
rect 7196 40562 7252 40572
rect 7308 40068 7364 41022
rect 7420 40852 7476 43486
rect 7532 43538 7588 43708
rect 7644 43650 7700 44492
rect 7868 44100 7924 44110
rect 7868 44006 7924 44044
rect 7644 43598 7646 43650
rect 7698 43598 7700 43650
rect 7644 43586 7700 43598
rect 7532 43486 7534 43538
rect 7586 43486 7588 43538
rect 7532 42868 7588 43486
rect 7644 42868 7700 42878
rect 7532 42866 7700 42868
rect 7532 42814 7646 42866
rect 7698 42814 7700 42866
rect 7532 42812 7700 42814
rect 7644 42802 7700 42812
rect 7420 40786 7476 40796
rect 7868 42754 7924 42766
rect 7868 42702 7870 42754
rect 7922 42702 7924 42754
rect 7532 40516 7588 40526
rect 7532 40422 7588 40460
rect 7308 40002 7364 40012
rect 7308 39620 7364 39630
rect 7364 39564 7700 39620
rect 7308 39526 7364 39564
rect 6860 39454 6862 39506
rect 6914 39454 6916 39506
rect 6860 39442 6916 39454
rect 7532 39396 7588 39406
rect 7532 39302 7588 39340
rect 7644 38946 7700 39564
rect 7644 38894 7646 38946
rect 7698 38894 7700 38946
rect 6972 37492 7028 37502
rect 7644 37492 7700 38894
rect 7868 39172 7924 42702
rect 7980 41858 8036 48188
rect 8652 47460 8708 52220
rect 8764 52182 8820 52220
rect 9324 52164 9380 52174
rect 9324 52070 9380 52108
rect 9548 51380 9604 53678
rect 9996 53732 10052 53742
rect 9996 53730 10724 53732
rect 9996 53678 9998 53730
rect 10050 53678 10724 53730
rect 9996 53676 10724 53678
rect 9996 53666 10052 53676
rect 10668 53508 10724 53676
rect 11452 53620 11508 54348
rect 11900 54310 11956 54348
rect 11900 53620 11956 53630
rect 11452 53618 11956 53620
rect 11452 53566 11902 53618
rect 11954 53566 11956 53618
rect 11452 53564 11956 53566
rect 9772 53284 9828 53294
rect 9772 52274 9828 53228
rect 9772 52222 9774 52274
rect 9826 52222 9828 52274
rect 9772 52210 9828 52222
rect 10332 52946 10388 52958
rect 10332 52894 10334 52946
rect 10386 52894 10388 52946
rect 10332 52164 10388 52894
rect 10668 52274 10724 53452
rect 10892 53508 10948 53518
rect 11340 53508 11396 53518
rect 10892 53506 11396 53508
rect 10892 53454 10894 53506
rect 10946 53454 11342 53506
rect 11394 53454 11396 53506
rect 10892 53452 11396 53454
rect 10892 53396 10948 53452
rect 10892 53330 10948 53340
rect 11340 52948 11396 53452
rect 11900 53396 11956 53564
rect 11900 53330 11956 53340
rect 11340 52882 11396 52892
rect 11452 52834 11508 52846
rect 11452 52782 11454 52834
rect 11506 52782 11508 52834
rect 11116 52388 11172 52398
rect 11116 52294 11172 52332
rect 10668 52222 10670 52274
rect 10722 52222 10724 52274
rect 10668 52210 10724 52222
rect 10780 52276 10836 52286
rect 9996 51492 10052 51502
rect 9996 51398 10052 51436
rect 10332 51380 10388 52108
rect 9548 51314 9604 51324
rect 10108 51378 10388 51380
rect 10108 51326 10334 51378
rect 10386 51326 10388 51378
rect 10108 51324 10388 51326
rect 10108 51044 10164 51324
rect 10332 51314 10388 51324
rect 10444 52162 10500 52174
rect 10444 52110 10446 52162
rect 10498 52110 10500 52162
rect 9996 50988 10164 51044
rect 9548 50708 9604 50718
rect 9548 50614 9604 50652
rect 9100 50596 9156 50606
rect 9100 50594 9268 50596
rect 9100 50542 9102 50594
rect 9154 50542 9268 50594
rect 9100 50540 9268 50542
rect 9100 50530 9156 50540
rect 8764 50372 8820 50382
rect 8764 50370 9044 50372
rect 8764 50318 8766 50370
rect 8818 50318 9044 50370
rect 8764 50316 9044 50318
rect 8764 50306 8820 50316
rect 8876 49812 8932 49822
rect 8876 49718 8932 49756
rect 8988 49698 9044 50316
rect 8988 49646 8990 49698
rect 9042 49646 9044 49698
rect 8764 48804 8820 48814
rect 8764 48242 8820 48748
rect 8988 48580 9044 49646
rect 8764 48190 8766 48242
rect 8818 48190 8820 48242
rect 8764 48178 8820 48190
rect 8876 48524 9044 48580
rect 9212 49026 9268 50540
rect 9996 50428 10052 50988
rect 9772 50372 10052 50428
rect 10108 50484 10164 50494
rect 9548 49812 9604 49822
rect 9548 49718 9604 49756
rect 9212 48974 9214 49026
rect 9266 48974 9268 49026
rect 8652 47404 8820 47460
rect 8652 47236 8708 47246
rect 8540 46452 8596 46462
rect 8540 46358 8596 46396
rect 8092 45890 8148 45902
rect 8092 45838 8094 45890
rect 8146 45838 8148 45890
rect 8092 45556 8148 45838
rect 8092 45490 8148 45500
rect 8652 44436 8708 47180
rect 8764 46786 8820 47404
rect 8876 47236 8932 48524
rect 8876 47170 8932 47180
rect 8988 48356 9044 48366
rect 9212 48356 9268 48974
rect 9548 49026 9604 49038
rect 9548 48974 9550 49026
rect 9602 48974 9604 49026
rect 9548 48804 9604 48974
rect 9772 49026 9828 50372
rect 10108 50260 10164 50428
rect 10444 50484 10500 52110
rect 10780 52162 10836 52220
rect 10780 52110 10782 52162
rect 10834 52110 10836 52162
rect 10780 52098 10836 52110
rect 11452 51716 11508 52782
rect 11228 51660 11452 51716
rect 11116 51380 11172 51390
rect 11116 51286 11172 51324
rect 10444 50418 10500 50428
rect 10668 51266 10724 51278
rect 10668 51214 10670 51266
rect 10722 51214 10724 51266
rect 9996 50204 10164 50260
rect 10332 50370 10388 50382
rect 10332 50318 10334 50370
rect 10386 50318 10388 50370
rect 9996 49698 10052 50204
rect 9996 49646 9998 49698
rect 10050 49646 10052 49698
rect 9996 49634 10052 49646
rect 10332 49700 10388 50318
rect 10332 49644 10612 49700
rect 10444 49476 10500 49486
rect 9772 48974 9774 49026
rect 9826 48974 9828 49026
rect 9772 48962 9828 48974
rect 9884 49250 9940 49262
rect 9884 49198 9886 49250
rect 9938 49198 9940 49250
rect 9548 48580 9604 48748
rect 9884 48580 9940 49198
rect 9548 48524 9828 48580
rect 8988 48354 9268 48356
rect 8988 48302 8990 48354
rect 9042 48302 9268 48354
rect 8988 48300 9268 48302
rect 8764 46734 8766 46786
rect 8818 46734 8820 46786
rect 8764 45780 8820 46734
rect 8876 46452 8932 46462
rect 8876 46358 8932 46396
rect 8876 45892 8932 45902
rect 8876 45798 8932 45836
rect 8764 45686 8820 45724
rect 8428 44380 8708 44436
rect 8092 43764 8148 43774
rect 8092 43670 8148 43708
rect 8204 43540 8260 43550
rect 8204 41972 8260 43484
rect 8316 42644 8372 42654
rect 8316 42550 8372 42588
rect 8204 41916 8372 41972
rect 7980 41806 7982 41858
rect 8034 41806 8036 41858
rect 7980 40852 8036 41806
rect 8204 41748 8260 41758
rect 8204 41654 8260 41692
rect 7980 40786 8036 40796
rect 8316 41186 8372 41916
rect 8316 41134 8318 41186
rect 8370 41134 8372 41186
rect 8204 40290 8260 40302
rect 8204 40238 8206 40290
rect 8258 40238 8260 40290
rect 8092 40180 8148 40190
rect 7980 39618 8036 39630
rect 7980 39566 7982 39618
rect 8034 39566 8036 39618
rect 7980 39284 8036 39566
rect 8092 39396 8148 40124
rect 8204 39620 8260 40238
rect 8204 39506 8260 39564
rect 8204 39454 8206 39506
rect 8258 39454 8260 39506
rect 8204 39442 8260 39454
rect 8092 39330 8148 39340
rect 7980 39218 8036 39228
rect 7868 38722 7924 39116
rect 7868 38670 7870 38722
rect 7922 38670 7924 38722
rect 7868 38658 7924 38670
rect 6972 37490 7700 37492
rect 6972 37438 6974 37490
rect 7026 37438 7646 37490
rect 7698 37438 7700 37490
rect 6972 37436 7700 37438
rect 8316 37940 8372 41134
rect 8428 41076 8484 44380
rect 8988 42308 9044 48300
rect 9548 47570 9604 47582
rect 9548 47518 9550 47570
rect 9602 47518 9604 47570
rect 9212 47234 9268 47246
rect 9212 47182 9214 47234
rect 9266 47182 9268 47234
rect 9212 46676 9268 47182
rect 9212 46610 9268 46620
rect 9548 45890 9604 47518
rect 9548 45838 9550 45890
rect 9602 45838 9604 45890
rect 9436 45668 9492 45678
rect 9436 45574 9492 45612
rect 9548 45444 9604 45838
rect 9548 45378 9604 45388
rect 9660 46676 9716 46686
rect 9548 43540 9604 43550
rect 9548 43446 9604 43484
rect 9212 42530 9268 42542
rect 9212 42478 9214 42530
rect 9266 42478 9268 42530
rect 9212 42308 9268 42478
rect 8876 42252 9268 42308
rect 8540 42196 8596 42206
rect 8540 42102 8596 42140
rect 8540 41300 8596 41310
rect 8876 41300 8932 42252
rect 8540 41298 8932 41300
rect 8540 41246 8542 41298
rect 8594 41246 8932 41298
rect 8540 41244 8932 41246
rect 8540 41234 8596 41244
rect 8988 41186 9044 41198
rect 8988 41134 8990 41186
rect 9042 41134 9044 41186
rect 8428 41020 8820 41076
rect 8428 40178 8484 40190
rect 8428 40126 8430 40178
rect 8482 40126 8484 40178
rect 8428 40068 8484 40126
rect 8484 40012 8708 40068
rect 8428 40002 8484 40012
rect 8652 39618 8708 40012
rect 8652 39566 8654 39618
rect 8706 39566 8708 39618
rect 8652 39554 8708 39566
rect 8428 39284 8484 39294
rect 8428 38722 8484 39228
rect 8428 38670 8430 38722
rect 8482 38670 8484 38722
rect 8428 38668 8484 38670
rect 8764 38668 8820 41020
rect 8876 40740 8932 40750
rect 8876 40626 8932 40684
rect 8876 40574 8878 40626
rect 8930 40574 8932 40626
rect 8876 40562 8932 40574
rect 8988 40292 9044 41134
rect 8988 40226 9044 40236
rect 9212 41074 9268 41086
rect 9212 41022 9214 41074
rect 9266 41022 9268 41074
rect 9212 40180 9268 41022
rect 9660 41074 9716 46620
rect 9772 46674 9828 48524
rect 9884 48514 9940 48524
rect 9772 46622 9774 46674
rect 9826 46622 9828 46674
rect 9772 44324 9828 46622
rect 9884 48242 9940 48254
rect 9884 48190 9886 48242
rect 9938 48190 9940 48242
rect 9884 45892 9940 48190
rect 10444 48242 10500 49420
rect 10556 49252 10612 49644
rect 10556 49138 10612 49196
rect 10556 49086 10558 49138
rect 10610 49086 10612 49138
rect 10556 49074 10612 49086
rect 10668 48356 10724 51214
rect 10668 48290 10724 48300
rect 10780 50370 10836 50382
rect 10780 50318 10782 50370
rect 10834 50318 10836 50370
rect 10444 48190 10446 48242
rect 10498 48190 10500 48242
rect 10444 48178 10500 48190
rect 10780 48132 10836 50318
rect 11116 50370 11172 50382
rect 11116 50318 11118 50370
rect 11170 50318 11172 50370
rect 11004 49810 11060 49822
rect 11004 49758 11006 49810
rect 11058 49758 11060 49810
rect 11004 49138 11060 49758
rect 11116 49252 11172 50318
rect 11116 49186 11172 49196
rect 11004 49086 11006 49138
rect 11058 49086 11060 49138
rect 11004 49074 11060 49086
rect 10892 48914 10948 48926
rect 10892 48862 10894 48914
rect 10946 48862 10948 48914
rect 10892 48468 10948 48862
rect 11116 48804 11172 48814
rect 11116 48710 11172 48748
rect 10892 48402 10948 48412
rect 11228 48244 11284 51660
rect 11452 51650 11508 51660
rect 11676 50370 11732 50382
rect 12012 50372 12068 54684
rect 12460 54628 12516 55020
rect 12460 54562 12516 54572
rect 12460 54404 12516 54414
rect 12348 54402 12516 54404
rect 12348 54350 12462 54402
rect 12514 54350 12516 54402
rect 12348 54348 12516 54350
rect 12236 53618 12292 53630
rect 12236 53566 12238 53618
rect 12290 53566 12292 53618
rect 12124 52948 12180 52958
rect 12124 52052 12180 52892
rect 12236 52500 12292 53566
rect 12348 52724 12404 54348
rect 12460 54338 12516 54348
rect 12348 52658 12404 52668
rect 12460 53844 12516 53854
rect 12572 53844 12628 56028
rect 12908 55972 12964 55982
rect 12460 53842 12628 53844
rect 12460 53790 12462 53842
rect 12514 53790 12628 53842
rect 12460 53788 12628 53790
rect 12796 55748 12852 55758
rect 12348 52500 12404 52510
rect 12236 52444 12348 52500
rect 12348 52274 12404 52444
rect 12460 52388 12516 53788
rect 12796 53730 12852 55692
rect 12908 55074 12964 55916
rect 14140 55972 14196 55982
rect 14140 55878 14196 55916
rect 14700 55970 14756 55982
rect 14700 55918 14702 55970
rect 14754 55918 14756 55970
rect 14700 55468 14756 55918
rect 14140 55412 14196 55422
rect 14140 55318 14196 55356
rect 14588 55412 14756 55468
rect 15036 55412 15092 57708
rect 25004 57540 25060 57550
rect 22988 57428 23044 57438
rect 22876 57372 22988 57428
rect 21084 57316 21140 57326
rect 16380 57204 16436 57214
rect 15596 56196 15652 56206
rect 15148 55970 15204 55982
rect 15148 55918 15150 55970
rect 15202 55918 15204 55970
rect 15148 55860 15204 55918
rect 15596 55970 15652 56140
rect 15596 55918 15598 55970
rect 15650 55918 15652 55970
rect 15148 55858 15316 55860
rect 15148 55806 15150 55858
rect 15202 55806 15316 55858
rect 15148 55804 15316 55806
rect 15148 55794 15204 55804
rect 15260 55412 15316 55804
rect 14588 55300 14644 55412
rect 15036 55356 15204 55412
rect 14588 55234 14644 55244
rect 14924 55300 14980 55310
rect 14980 55244 15092 55300
rect 14924 55234 14980 55244
rect 15036 55186 15092 55244
rect 15036 55134 15038 55186
rect 15090 55134 15092 55186
rect 15036 55122 15092 55134
rect 12908 55022 12910 55074
rect 12962 55022 12964 55074
rect 12908 54740 12964 55022
rect 13916 55074 13972 55086
rect 13916 55022 13918 55074
rect 13970 55022 13972 55074
rect 13916 54740 13972 55022
rect 14700 55076 14756 55086
rect 14700 55074 14980 55076
rect 14700 55022 14702 55074
rect 14754 55022 14980 55074
rect 14700 55020 14980 55022
rect 13916 54684 14420 54740
rect 12908 54674 12964 54684
rect 13692 54516 13748 54526
rect 14028 54516 14084 54526
rect 14252 54516 14308 54526
rect 13692 54514 14252 54516
rect 13692 54462 13694 54514
rect 13746 54462 14030 54514
rect 14082 54462 14252 54514
rect 13692 54460 14252 54462
rect 13692 54450 13748 54460
rect 14028 54450 14084 54460
rect 14252 54450 14308 54460
rect 12908 54402 12964 54414
rect 12908 54350 12910 54402
rect 12962 54350 12964 54402
rect 12908 54068 12964 54350
rect 12908 54002 12964 54012
rect 13356 54402 13412 54414
rect 13356 54350 13358 54402
rect 13410 54350 13412 54402
rect 12796 53678 12798 53730
rect 12850 53678 12852 53730
rect 12796 53666 12852 53678
rect 13132 53956 13188 53966
rect 12572 52948 12628 52958
rect 12572 52854 12628 52892
rect 12460 52322 12516 52332
rect 12348 52222 12350 52274
rect 12402 52222 12404 52274
rect 12348 52210 12404 52222
rect 12572 52164 12628 52174
rect 12572 52162 12740 52164
rect 12572 52110 12574 52162
rect 12626 52110 12740 52162
rect 12572 52108 12740 52110
rect 12572 52098 12628 52108
rect 12460 52052 12516 52062
rect 12124 52050 12516 52052
rect 12124 51998 12462 52050
rect 12514 51998 12516 52050
rect 12124 51996 12516 51998
rect 12348 51716 12404 51726
rect 12236 51266 12292 51278
rect 12236 51214 12238 51266
rect 12290 51214 12292 51266
rect 12236 50596 12292 51214
rect 12348 50708 12404 51660
rect 12460 51156 12516 51996
rect 12684 51380 12740 52108
rect 12684 51286 12740 51324
rect 12460 51100 12740 51156
rect 12460 50708 12516 50718
rect 12348 50706 12516 50708
rect 12348 50654 12462 50706
rect 12514 50654 12516 50706
rect 12348 50652 12516 50654
rect 12460 50642 12516 50652
rect 12236 50530 12292 50540
rect 11676 50318 11678 50370
rect 11730 50318 11732 50370
rect 11676 50148 11732 50318
rect 11676 50082 11732 50092
rect 11900 50370 12068 50372
rect 11900 50318 12014 50370
rect 12066 50318 12068 50370
rect 11900 50316 12068 50318
rect 11340 49810 11396 49822
rect 11340 49758 11342 49810
rect 11394 49758 11396 49810
rect 11340 48468 11396 49758
rect 11452 49698 11508 49710
rect 11452 49646 11454 49698
rect 11506 49646 11508 49698
rect 11452 49364 11508 49646
rect 11452 49298 11508 49308
rect 11564 49028 11620 49038
rect 11788 49028 11844 49038
rect 11340 48412 11508 48468
rect 10556 48076 10836 48132
rect 11004 48242 11284 48244
rect 11004 48190 11230 48242
rect 11282 48190 11284 48242
rect 11004 48188 11284 48190
rect 9996 47236 10052 47246
rect 9996 47142 10052 47180
rect 10556 47012 10612 48076
rect 11004 47908 11060 48188
rect 11228 48178 11284 48188
rect 11340 48242 11396 48254
rect 11340 48190 11342 48242
rect 11394 48190 11396 48242
rect 10668 47852 11060 47908
rect 10668 47570 10724 47852
rect 10668 47518 10670 47570
rect 10722 47518 10724 47570
rect 10668 47506 10724 47518
rect 11004 47460 11060 47470
rect 11004 47458 11284 47460
rect 11004 47406 11006 47458
rect 11058 47406 11284 47458
rect 11004 47404 11284 47406
rect 11004 47394 11060 47404
rect 10556 46956 10724 47012
rect 9884 45826 9940 45836
rect 9996 46786 10052 46798
rect 9996 46734 9998 46786
rect 10050 46734 10052 46786
rect 9996 45108 10052 46734
rect 10556 46786 10612 46798
rect 10556 46734 10558 46786
rect 10610 46734 10612 46786
rect 10332 46676 10388 46686
rect 10332 46582 10388 46620
rect 10332 46002 10388 46014
rect 10332 45950 10334 46002
rect 10386 45950 10388 46002
rect 9996 45042 10052 45052
rect 10108 45890 10164 45902
rect 10108 45838 10110 45890
rect 10162 45838 10164 45890
rect 10108 45106 10164 45838
rect 10108 45054 10110 45106
rect 10162 45054 10164 45106
rect 9996 44324 10052 44334
rect 9772 44322 10052 44324
rect 9772 44270 9998 44322
rect 10050 44270 10052 44322
rect 9772 44268 10052 44270
rect 9996 44258 10052 44268
rect 10108 44098 10164 45054
rect 10332 44324 10388 45950
rect 10444 45892 10500 45902
rect 10444 45778 10500 45836
rect 10444 45726 10446 45778
rect 10498 45726 10500 45778
rect 10444 45218 10500 45726
rect 10444 45166 10446 45218
rect 10498 45166 10500 45218
rect 10444 45154 10500 45166
rect 10332 44268 10500 44324
rect 10108 44046 10110 44098
rect 10162 44046 10164 44098
rect 10108 43428 10164 44046
rect 10332 44098 10388 44110
rect 10332 44046 10334 44098
rect 10386 44046 10388 44098
rect 10332 43988 10388 44046
rect 10332 43922 10388 43932
rect 10332 43428 10388 43438
rect 10108 43426 10388 43428
rect 10108 43374 10334 43426
rect 10386 43374 10388 43426
rect 10108 43372 10388 43374
rect 10332 42754 10388 43372
rect 10332 42702 10334 42754
rect 10386 42702 10388 42754
rect 10332 42690 10388 42702
rect 9772 42642 9828 42654
rect 9772 42590 9774 42642
rect 9826 42590 9828 42642
rect 9772 41188 9828 42590
rect 9772 41122 9828 41132
rect 10332 41972 10388 41982
rect 9660 41022 9662 41074
rect 9714 41022 9716 41074
rect 9660 40852 9716 41022
rect 9660 40786 9716 40796
rect 9772 40964 9828 40974
rect 9212 39618 9268 40124
rect 9772 39842 9828 40908
rect 9884 40628 9940 40638
rect 9884 40534 9940 40572
rect 10220 40516 10276 40526
rect 10108 40404 10164 40414
rect 10108 40310 10164 40348
rect 9772 39790 9774 39842
rect 9826 39790 9828 39842
rect 9772 39778 9828 39790
rect 9212 39566 9214 39618
rect 9266 39566 9268 39618
rect 9212 39060 9268 39566
rect 9996 39620 10052 39630
rect 9996 39526 10052 39564
rect 9548 39060 9604 39070
rect 9212 39058 9604 39060
rect 9212 39006 9550 39058
rect 9602 39006 9604 39058
rect 9212 39004 9604 39006
rect 9548 38994 9604 39004
rect 8428 38612 8820 38668
rect 9996 38948 10052 38958
rect 9996 38722 10052 38892
rect 9996 38670 9998 38722
rect 10050 38670 10052 38722
rect 9996 38658 10052 38670
rect 10220 38668 10276 40460
rect 10332 39172 10388 41916
rect 10332 39106 10388 39116
rect 10220 38612 10388 38668
rect 8316 37492 8372 37884
rect 8652 37492 8708 37502
rect 8316 37490 8708 37492
rect 8316 37438 8654 37490
rect 8706 37438 8708 37490
rect 8316 37436 8708 37438
rect 6972 37426 7028 37436
rect 7644 37426 7700 37436
rect 8652 37426 8708 37436
rect 7196 37268 7252 37278
rect 7196 37174 7252 37212
rect 8428 37268 8484 37278
rect 6412 36866 6468 36876
rect 8204 37154 8260 37166
rect 8204 37102 8206 37154
rect 8258 37102 8260 37154
rect 8204 36484 8260 37102
rect 8204 36418 8260 36428
rect 8428 36482 8484 37212
rect 8428 36430 8430 36482
rect 8482 36430 8484 36482
rect 8428 36418 8484 36430
rect 7532 36370 7588 36382
rect 7532 36318 7534 36370
rect 7586 36318 7588 36370
rect 7420 36148 7476 36158
rect 6860 35698 6916 35710
rect 6860 35646 6862 35698
rect 6914 35646 6916 35698
rect 6860 35588 6916 35646
rect 7420 35698 7476 36092
rect 7420 35646 7422 35698
rect 7474 35646 7476 35698
rect 7420 35634 7476 35646
rect 6860 35522 6916 35532
rect 6300 34692 6356 34702
rect 6300 34598 6356 34636
rect 5628 34402 5684 34412
rect 6076 34244 6132 34254
rect 4844 34132 4900 34142
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 1708 33234 1764 33246
rect 1708 33182 1710 33234
rect 1762 33182 1764 33234
rect 1708 33012 1764 33182
rect 2044 33236 2100 33246
rect 2044 33142 2100 33180
rect 1708 32946 1764 32956
rect 2492 33122 2548 33134
rect 2492 33070 2494 33122
rect 2546 33070 2548 33122
rect 2492 33012 2548 33070
rect 2492 32946 2548 32956
rect 1820 32450 1876 32462
rect 1820 32398 1822 32450
rect 1874 32398 1876 32450
rect 1820 31778 1876 32398
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 1820 31726 1822 31778
rect 1874 31726 1876 31778
rect 1820 30996 1876 31726
rect 2380 31668 2436 31678
rect 2380 31574 2436 31612
rect 2044 31556 2100 31566
rect 2044 31462 2100 31500
rect 4620 31554 4676 31566
rect 4620 31502 4622 31554
rect 4674 31502 4676 31554
rect 1820 30930 1876 30940
rect 4284 30996 4340 31006
rect 4620 30996 4676 31502
rect 4284 30994 4676 30996
rect 4284 30942 4286 30994
rect 4338 30942 4676 30994
rect 4284 30940 4676 30942
rect 4844 30994 4900 34076
rect 5516 34132 5572 34142
rect 5516 34038 5572 34076
rect 6076 34130 6132 34188
rect 6076 34078 6078 34130
rect 6130 34078 6132 34130
rect 6076 34066 6132 34078
rect 6636 33908 6692 33918
rect 4844 30942 4846 30994
rect 4898 30942 4900 30994
rect 1932 30770 1988 30782
rect 1932 30718 1934 30770
rect 1986 30718 1988 30770
rect 1932 30324 1988 30718
rect 4284 30772 4340 30940
rect 4284 30706 4340 30716
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 1932 30258 1988 30268
rect 4172 30210 4228 30222
rect 4172 30158 4174 30210
rect 4226 30158 4228 30210
rect 2492 30098 2548 30110
rect 2492 30046 2494 30098
rect 2546 30046 2548 30098
rect 2492 29652 2548 30046
rect 2492 29586 2548 29596
rect 1932 29204 1988 29214
rect 1932 29110 1988 29148
rect 1932 28754 1988 28766
rect 1932 28702 1934 28754
rect 1986 28702 1988 28754
rect 1932 28308 1988 28702
rect 4172 28532 4228 30158
rect 4284 29426 4340 29438
rect 4284 29374 4286 29426
rect 4338 29374 4340 29426
rect 4284 28868 4340 29374
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4284 28802 4340 28812
rect 4284 28644 4340 28654
rect 4284 28550 4340 28588
rect 4172 28466 4228 28476
rect 1932 28242 1988 28252
rect 4620 27860 4676 27870
rect 4844 27860 4900 30942
rect 5404 30996 5460 31006
rect 6636 30996 6692 33852
rect 7532 33236 7588 36318
rect 7868 36260 7924 36270
rect 7868 36166 7924 36204
rect 8204 35924 8260 35934
rect 8092 35922 8260 35924
rect 8092 35870 8206 35922
rect 8258 35870 8260 35922
rect 8092 35868 8260 35870
rect 7532 33170 7588 33180
rect 7868 34692 7924 34702
rect 5404 30994 5684 30996
rect 5404 30942 5406 30994
rect 5458 30942 5684 30994
rect 5404 30940 5684 30942
rect 5404 30930 5460 30940
rect 5628 30098 5684 30940
rect 6636 30930 6692 30940
rect 7868 31218 7924 34636
rect 8092 34020 8148 35868
rect 8204 35858 8260 35868
rect 8428 35698 8484 35710
rect 8428 35646 8430 35698
rect 8482 35646 8484 35698
rect 8428 34804 8484 35646
rect 8428 34738 8484 34748
rect 8540 35364 8596 35374
rect 8316 34692 8372 34702
rect 8316 34356 8372 34636
rect 8316 34262 8372 34300
rect 8092 33954 8148 33964
rect 8316 34132 8372 34142
rect 8316 33460 8372 34076
rect 8316 33458 8484 33460
rect 8316 33406 8318 33458
rect 8370 33406 8484 33458
rect 8316 33404 8484 33406
rect 8316 33394 8372 33404
rect 8428 32228 8484 33404
rect 8540 33234 8596 35308
rect 8764 35028 8820 38612
rect 10220 37940 10276 37950
rect 10220 37846 10276 37884
rect 8876 37266 8932 37278
rect 8876 37214 8878 37266
rect 8930 37214 8932 37266
rect 8876 35700 8932 37214
rect 9660 37266 9716 37278
rect 9660 37214 9662 37266
rect 9714 37214 9716 37266
rect 8988 36596 9044 36606
rect 8988 36502 9044 36540
rect 9436 36482 9492 36494
rect 9436 36430 9438 36482
rect 9490 36430 9492 36482
rect 8988 35700 9044 35710
rect 8876 35644 8988 35700
rect 8988 35634 9044 35644
rect 9436 35364 9492 36430
rect 9436 35298 9492 35308
rect 9660 36484 9716 37214
rect 9996 37268 10052 37278
rect 10332 37268 10388 38612
rect 10444 37604 10500 44268
rect 10556 41412 10612 46734
rect 10668 42756 10724 46956
rect 11228 46786 11284 47404
rect 11340 47124 11396 48190
rect 11452 47796 11508 48412
rect 11564 48466 11620 48972
rect 11564 48414 11566 48466
rect 11618 48414 11620 48466
rect 11564 48402 11620 48414
rect 11676 49026 11844 49028
rect 11676 48974 11790 49026
rect 11842 48974 11844 49026
rect 11676 48972 11844 48974
rect 11452 47730 11508 47740
rect 11564 48132 11620 48142
rect 11676 48132 11732 48972
rect 11788 48962 11844 48972
rect 11564 48130 11732 48132
rect 11564 48078 11566 48130
rect 11618 48078 11732 48130
rect 11564 48076 11732 48078
rect 11452 47572 11508 47582
rect 11452 47478 11508 47516
rect 11452 47124 11508 47134
rect 11340 47068 11452 47124
rect 11452 47058 11508 47068
rect 11564 46788 11620 48076
rect 11676 47684 11732 47694
rect 11676 46898 11732 47628
rect 11900 47068 11956 50316
rect 12012 50306 12068 50316
rect 12348 49810 12404 49822
rect 12348 49758 12350 49810
rect 12402 49758 12404 49810
rect 12012 49698 12068 49710
rect 12012 49646 12014 49698
rect 12066 49646 12068 49698
rect 12012 49476 12068 49646
rect 12012 49410 12068 49420
rect 12236 49028 12292 49038
rect 12348 49028 12404 49758
rect 12236 49026 12404 49028
rect 12236 48974 12238 49026
rect 12290 48974 12404 49026
rect 12236 48972 12404 48974
rect 12572 49252 12628 49262
rect 12572 49026 12628 49196
rect 12572 48974 12574 49026
rect 12626 48974 12628 49026
rect 12236 48804 12292 48972
rect 11676 46846 11678 46898
rect 11730 46846 11732 46898
rect 11676 46834 11732 46846
rect 11788 47012 11956 47068
rect 12012 47234 12068 47246
rect 12012 47182 12014 47234
rect 12066 47182 12068 47234
rect 11228 46734 11230 46786
rect 11282 46734 11284 46786
rect 11228 45332 11284 46734
rect 11228 45266 11284 45276
rect 11452 46732 11620 46788
rect 11228 43988 11284 43998
rect 11116 43540 11172 43550
rect 10668 42690 10724 42700
rect 11004 43538 11172 43540
rect 11004 43486 11118 43538
rect 11170 43486 11172 43538
rect 11004 43484 11172 43486
rect 10892 42642 10948 42654
rect 10892 42590 10894 42642
rect 10946 42590 10948 42642
rect 10780 42082 10836 42094
rect 10780 42030 10782 42082
rect 10834 42030 10836 42082
rect 10668 41972 10724 41982
rect 10780 41972 10836 42030
rect 10724 41916 10836 41972
rect 10668 41906 10724 41916
rect 10556 41356 10836 41412
rect 10556 41186 10612 41198
rect 10556 41134 10558 41186
rect 10610 41134 10612 41186
rect 10556 40964 10612 41134
rect 10556 40898 10612 40908
rect 10668 40292 10724 40302
rect 10668 39732 10724 40236
rect 10668 39618 10724 39676
rect 10668 39566 10670 39618
rect 10722 39566 10724 39618
rect 10668 39554 10724 39566
rect 10780 39058 10836 41356
rect 10892 40516 10948 42590
rect 11004 40964 11060 43484
rect 11116 43474 11172 43484
rect 11116 43314 11172 43326
rect 11116 43262 11118 43314
rect 11170 43262 11172 43314
rect 11116 41748 11172 43262
rect 11116 41682 11172 41692
rect 11004 40898 11060 40908
rect 10892 40450 10948 40460
rect 10780 39006 10782 39058
rect 10834 39006 10836 39058
rect 10556 37828 10612 37838
rect 10556 37734 10612 37772
rect 10444 37538 10500 37548
rect 10668 37268 10724 37278
rect 10332 37212 10668 37268
rect 9996 37154 10052 37212
rect 10668 37174 10724 37212
rect 9996 37102 9998 37154
rect 10050 37102 10052 37154
rect 9772 36484 9828 36494
rect 9660 36482 9828 36484
rect 9660 36430 9774 36482
rect 9826 36430 9828 36482
rect 9660 36428 9828 36430
rect 8764 34962 8820 34972
rect 8652 34916 8708 34926
rect 8652 34822 8708 34860
rect 8988 34914 9044 34926
rect 8988 34862 8990 34914
rect 9042 34862 9044 34914
rect 8988 34692 9044 34862
rect 9436 34804 9492 34814
rect 9436 34710 9492 34748
rect 8988 34132 9044 34636
rect 9100 34356 9156 34366
rect 9660 34356 9716 36428
rect 9772 36418 9828 36428
rect 9996 35698 10052 37102
rect 10444 36260 10500 36270
rect 9996 35646 9998 35698
rect 10050 35646 10052 35698
rect 9996 35634 10052 35646
rect 10108 35700 10164 35710
rect 10108 35586 10164 35644
rect 10108 35534 10110 35586
rect 10162 35534 10164 35586
rect 10108 35522 10164 35534
rect 10444 34802 10500 36204
rect 10668 35812 10724 35822
rect 10780 35812 10836 39006
rect 11228 38724 11284 43932
rect 11452 43314 11508 46732
rect 11564 46564 11620 46574
rect 11788 46564 11844 47012
rect 11564 46562 11844 46564
rect 11564 46510 11566 46562
rect 11618 46510 11844 46562
rect 11564 46508 11844 46510
rect 11900 46786 11956 46798
rect 11900 46734 11902 46786
rect 11954 46734 11956 46786
rect 11900 46564 11956 46734
rect 12012 46676 12068 47182
rect 12012 46582 12068 46620
rect 11564 46116 11620 46508
rect 11564 46050 11620 46060
rect 11676 45892 11732 45902
rect 11676 45218 11732 45836
rect 11788 45890 11844 45902
rect 11788 45838 11790 45890
rect 11842 45838 11844 45890
rect 11788 45780 11844 45838
rect 11788 45714 11844 45724
rect 11676 45166 11678 45218
rect 11730 45166 11732 45218
rect 11676 45154 11732 45166
rect 11788 45332 11844 45342
rect 11788 45106 11844 45276
rect 11788 45054 11790 45106
rect 11842 45054 11844 45106
rect 11788 45042 11844 45054
rect 11452 43262 11454 43314
rect 11506 43262 11508 43314
rect 11452 42196 11508 43262
rect 11788 44436 11844 44446
rect 11452 42130 11508 42140
rect 11564 42756 11620 42766
rect 11340 41972 11396 41982
rect 11340 41878 11396 41916
rect 11452 41186 11508 41198
rect 11452 41134 11454 41186
rect 11506 41134 11508 41186
rect 11340 41076 11396 41086
rect 11340 40402 11396 41020
rect 11340 40350 11342 40402
rect 11394 40350 11396 40402
rect 11340 39842 11396 40350
rect 11452 40404 11508 41134
rect 11452 40338 11508 40348
rect 11340 39790 11342 39842
rect 11394 39790 11396 39842
rect 11340 39778 11396 39790
rect 11564 39396 11620 42700
rect 11676 42308 11732 42318
rect 11676 41298 11732 42252
rect 11676 41246 11678 41298
rect 11730 41246 11732 41298
rect 11676 41234 11732 41246
rect 11340 38836 11396 38846
rect 11564 38836 11620 39340
rect 11340 38834 11620 38836
rect 11340 38782 11342 38834
rect 11394 38782 11620 38834
rect 11340 38780 11620 38782
rect 11676 40404 11732 40414
rect 11676 39058 11732 40348
rect 11676 39006 11678 39058
rect 11730 39006 11732 39058
rect 11340 38770 11396 38780
rect 11676 38668 11732 39006
rect 11228 38658 11284 38668
rect 11340 38612 11732 38668
rect 11340 37492 11396 38612
rect 11004 37436 11396 37492
rect 11004 36594 11060 37436
rect 11004 36542 11006 36594
rect 11058 36542 11060 36594
rect 11004 36530 11060 36542
rect 11116 37266 11172 37278
rect 11116 37214 11118 37266
rect 11170 37214 11172 37266
rect 11116 36148 11172 37214
rect 11788 36596 11844 44380
rect 11900 43988 11956 46508
rect 12236 45332 12292 48748
rect 12348 48580 12404 48590
rect 12348 48244 12404 48524
rect 12348 47458 12404 48188
rect 12460 48356 12516 48366
rect 12460 48242 12516 48300
rect 12460 48190 12462 48242
rect 12514 48190 12516 48242
rect 12460 48178 12516 48190
rect 12348 47406 12350 47458
rect 12402 47406 12404 47458
rect 12348 47394 12404 47406
rect 12460 46676 12516 46686
rect 12348 46674 12516 46676
rect 12348 46622 12462 46674
rect 12514 46622 12516 46674
rect 12348 46620 12516 46622
rect 12348 46564 12404 46620
rect 12460 46610 12516 46620
rect 12348 46498 12404 46508
rect 12236 45276 12516 45332
rect 11900 43922 11956 43932
rect 12348 44098 12404 44110
rect 12348 44046 12350 44098
rect 12402 44046 12404 44098
rect 12348 43540 12404 44046
rect 12124 43538 12404 43540
rect 12124 43486 12350 43538
rect 12402 43486 12404 43538
rect 12124 43484 12404 43486
rect 12124 42866 12180 43484
rect 12348 43474 12404 43484
rect 12460 43316 12516 45276
rect 12572 44100 12628 48974
rect 12684 44436 12740 51100
rect 13020 50370 13076 50382
rect 13020 50318 13022 50370
rect 13074 50318 13076 50370
rect 13020 50260 13076 50318
rect 13020 50194 13076 50204
rect 13020 49028 13076 49038
rect 13132 49028 13188 53900
rect 13356 53620 13412 54350
rect 13580 54404 13636 54414
rect 13580 54310 13636 54348
rect 13916 53732 13972 53742
rect 13356 53554 13412 53564
rect 13804 53730 13972 53732
rect 13804 53678 13918 53730
rect 13970 53678 13972 53730
rect 13804 53676 13972 53678
rect 13692 53506 13748 53518
rect 13692 53454 13694 53506
rect 13746 53454 13748 53506
rect 13692 53284 13748 53454
rect 13692 53218 13748 53228
rect 13356 53172 13412 53182
rect 13356 53078 13412 53116
rect 13804 53060 13860 53676
rect 13916 53666 13972 53676
rect 13692 53004 13860 53060
rect 13468 52386 13524 52398
rect 13468 52334 13470 52386
rect 13522 52334 13524 52386
rect 13244 51380 13300 51390
rect 13244 51266 13300 51324
rect 13244 51214 13246 51266
rect 13298 51214 13300 51266
rect 13244 51202 13300 51214
rect 13356 49924 13412 49934
rect 13020 49026 13188 49028
rect 13020 48974 13022 49026
rect 13074 48974 13188 49026
rect 13020 48972 13188 48974
rect 13244 49922 13412 49924
rect 13244 49870 13358 49922
rect 13410 49870 13412 49922
rect 13244 49868 13412 49870
rect 13020 48962 13076 48972
rect 12908 47458 12964 47470
rect 12908 47406 12910 47458
rect 12962 47406 12964 47458
rect 12908 46004 12964 47406
rect 13132 47460 13188 47470
rect 12908 45938 12964 45948
rect 13020 47012 13076 47022
rect 12908 45668 12964 45678
rect 13020 45668 13076 46956
rect 13132 46898 13188 47404
rect 13132 46846 13134 46898
rect 13186 46846 13188 46898
rect 13132 46834 13188 46846
rect 12908 45666 13076 45668
rect 12908 45614 12910 45666
rect 12962 45614 13076 45666
rect 12908 45612 13076 45614
rect 12908 45602 12964 45612
rect 12684 44370 12740 44380
rect 12908 45106 12964 45118
rect 12908 45054 12910 45106
rect 12962 45054 12964 45106
rect 12908 44324 12964 45054
rect 13020 45106 13076 45612
rect 13244 45556 13300 49868
rect 13356 49858 13412 49868
rect 13468 48692 13524 52334
rect 13580 50820 13636 50830
rect 13692 50820 13748 53004
rect 13916 52948 13972 52958
rect 13804 52836 13860 52846
rect 13804 52742 13860 52780
rect 13804 52386 13860 52398
rect 13804 52334 13806 52386
rect 13858 52334 13860 52386
rect 13804 52274 13860 52334
rect 13804 52222 13806 52274
rect 13858 52222 13860 52274
rect 13804 52210 13860 52222
rect 13916 51490 13972 52892
rect 14252 52948 14308 52958
rect 14252 52854 14308 52892
rect 14140 52834 14196 52846
rect 14140 52782 14142 52834
rect 14194 52782 14196 52834
rect 13916 51438 13918 51490
rect 13970 51438 13972 51490
rect 13692 50764 13860 50820
rect 13580 50706 13636 50764
rect 13580 50654 13582 50706
rect 13634 50654 13636 50706
rect 13580 49252 13636 50654
rect 13580 49186 13636 49196
rect 13692 50596 13748 50606
rect 13580 49028 13636 49038
rect 13580 48934 13636 48972
rect 13468 48636 13636 48692
rect 13468 48468 13524 48478
rect 13468 48242 13524 48412
rect 13468 48190 13470 48242
rect 13522 48190 13524 48242
rect 13468 48178 13524 48190
rect 13468 48018 13524 48030
rect 13468 47966 13470 48018
rect 13522 47966 13524 48018
rect 13468 47458 13524 47966
rect 13468 47406 13470 47458
rect 13522 47406 13524 47458
rect 13468 47394 13524 47406
rect 13580 47236 13636 48636
rect 13468 47180 13636 47236
rect 13356 47012 13412 47022
rect 13468 47012 13524 47180
rect 13412 46956 13524 47012
rect 13580 47012 13636 47022
rect 13356 46946 13412 46956
rect 13580 46898 13636 46956
rect 13580 46846 13582 46898
rect 13634 46846 13636 46898
rect 13580 46834 13636 46846
rect 13020 45054 13022 45106
rect 13074 45054 13076 45106
rect 13020 44996 13076 45054
rect 13020 44930 13076 44940
rect 13132 45500 13300 45556
rect 13468 45778 13524 45790
rect 13468 45726 13470 45778
rect 13522 45726 13524 45778
rect 13132 44660 13188 45500
rect 13244 45332 13300 45342
rect 13468 45332 13524 45726
rect 13244 45330 13524 45332
rect 13244 45278 13246 45330
rect 13298 45278 13524 45330
rect 13244 45276 13524 45278
rect 13244 45266 13300 45276
rect 13356 45108 13412 45118
rect 13356 45014 13412 45052
rect 13132 44604 13412 44660
rect 12908 44230 12964 44268
rect 12572 44044 12964 44100
rect 12124 42814 12126 42866
rect 12178 42814 12180 42866
rect 12124 41972 12180 42814
rect 12124 41878 12180 41916
rect 12348 43260 12516 43316
rect 12796 43876 12852 43886
rect 12012 40402 12068 40414
rect 12012 40350 12014 40402
rect 12066 40350 12068 40402
rect 11900 39620 11956 39630
rect 11900 39060 11956 39564
rect 11900 38994 11956 39004
rect 12012 38836 12068 40350
rect 12348 40404 12404 43260
rect 12684 42980 12740 42990
rect 12572 42868 12628 42878
rect 12572 42082 12628 42812
rect 12684 42866 12740 42924
rect 12684 42814 12686 42866
rect 12738 42814 12740 42866
rect 12684 42802 12740 42814
rect 12572 42030 12574 42082
rect 12626 42030 12628 42082
rect 12572 42018 12628 42030
rect 12460 41972 12516 41982
rect 12460 41878 12516 41916
rect 12684 41860 12740 41870
rect 12684 41186 12740 41804
rect 12684 41134 12686 41186
rect 12738 41134 12740 41186
rect 12684 41076 12740 41134
rect 12684 41010 12740 41020
rect 12796 40626 12852 43820
rect 12796 40574 12798 40626
rect 12850 40574 12852 40626
rect 12796 40562 12852 40574
rect 12684 40404 12740 40414
rect 12348 40402 12740 40404
rect 12348 40350 12686 40402
rect 12738 40350 12740 40402
rect 12348 40348 12740 40350
rect 12572 39060 12628 39070
rect 12572 38966 12628 39004
rect 12236 38836 12292 38846
rect 12012 38780 12236 38836
rect 12236 38742 12292 38780
rect 12684 37154 12740 40348
rect 12796 40292 12852 40302
rect 12796 39730 12852 40236
rect 12796 39678 12798 39730
rect 12850 39678 12852 39730
rect 12796 39666 12852 39678
rect 12908 39620 12964 44044
rect 13356 43538 13412 44604
rect 13580 44100 13636 44110
rect 13580 44006 13636 44044
rect 13356 43486 13358 43538
rect 13410 43486 13412 43538
rect 13356 41860 13412 43486
rect 13692 42756 13748 50540
rect 13804 50036 13860 50764
rect 13916 50428 13972 51438
rect 14028 52164 14084 52174
rect 14028 50820 14084 52108
rect 14140 51380 14196 52782
rect 14364 52276 14420 54684
rect 14476 54628 14532 54638
rect 14476 53730 14532 54572
rect 14700 54516 14756 55020
rect 14924 54738 14980 55020
rect 15148 54964 15204 55356
rect 14924 54686 14926 54738
rect 14978 54686 14980 54738
rect 14924 54674 14980 54686
rect 15036 54908 15204 54964
rect 14700 54450 14756 54460
rect 14476 53678 14478 53730
rect 14530 53678 14532 53730
rect 14476 53666 14532 53678
rect 14588 54402 14644 54414
rect 14588 54350 14590 54402
rect 14642 54350 14644 54402
rect 14364 52162 14420 52220
rect 14364 52110 14366 52162
rect 14418 52110 14420 52162
rect 14364 52098 14420 52110
rect 14476 53508 14532 53518
rect 14140 51314 14196 51324
rect 14252 51266 14308 51278
rect 14252 51214 14254 51266
rect 14306 51214 14308 51266
rect 14140 50820 14196 50830
rect 14028 50818 14196 50820
rect 14028 50766 14142 50818
rect 14194 50766 14196 50818
rect 14028 50764 14196 50766
rect 14140 50754 14196 50764
rect 14252 50708 14308 51214
rect 14476 51154 14532 53452
rect 14588 51492 14644 54350
rect 14812 53508 14868 53518
rect 14812 53414 14868 53452
rect 14588 51436 14868 51492
rect 14476 51102 14478 51154
rect 14530 51102 14532 51154
rect 14476 51090 14532 51102
rect 14252 50642 14308 50652
rect 13916 50372 14644 50428
rect 13804 49252 13860 49980
rect 14140 49810 14196 50372
rect 14588 50370 14644 50372
rect 14588 50318 14590 50370
rect 14642 50318 14644 50370
rect 14588 50306 14644 50318
rect 14140 49758 14142 49810
rect 14194 49758 14196 49810
rect 14140 49746 14196 49758
rect 14700 49698 14756 49710
rect 14700 49646 14702 49698
rect 14754 49646 14756 49698
rect 14700 49252 14756 49646
rect 13804 49196 14196 49252
rect 13916 49026 13972 49038
rect 13916 48974 13918 49026
rect 13970 48974 13972 49026
rect 13804 44884 13860 44894
rect 13804 44100 13860 44828
rect 13804 44034 13860 44044
rect 13916 43876 13972 48974
rect 14140 49028 14196 49196
rect 14700 49186 14756 49196
rect 14476 49028 14532 49038
rect 14140 49026 14532 49028
rect 14140 48974 14478 49026
rect 14530 48974 14532 49026
rect 14140 48972 14532 48974
rect 14028 48914 14084 48926
rect 14028 48862 14030 48914
rect 14082 48862 14084 48914
rect 14028 47346 14084 48862
rect 14028 47294 14030 47346
rect 14082 47294 14084 47346
rect 14028 47282 14084 47294
rect 14028 46788 14084 46798
rect 14028 46694 14084 46732
rect 14252 46452 14308 46462
rect 14364 46452 14420 48972
rect 14476 48962 14532 48972
rect 14588 49028 14644 49038
rect 14476 48356 14532 48366
rect 14476 47348 14532 48300
rect 14476 46786 14532 47292
rect 14476 46734 14478 46786
rect 14530 46734 14532 46786
rect 14476 46722 14532 46734
rect 14588 46786 14644 48972
rect 14812 48242 14868 51436
rect 15036 51380 15092 54908
rect 15260 51492 15316 55356
rect 15372 55300 15428 55310
rect 15372 55186 15428 55244
rect 15372 55134 15374 55186
rect 15426 55134 15428 55186
rect 15372 54628 15428 55134
rect 15596 55188 15652 55918
rect 16044 55970 16100 55982
rect 16044 55918 16046 55970
rect 16098 55918 16100 55970
rect 15932 55300 15988 55310
rect 15932 55206 15988 55244
rect 15596 55122 15652 55132
rect 15372 54562 15428 54572
rect 15484 54402 15540 54414
rect 15484 54350 15486 54402
rect 15538 54350 15540 54402
rect 15260 51426 15316 51436
rect 15372 53730 15428 53742
rect 15372 53678 15374 53730
rect 15426 53678 15428 53730
rect 14812 48190 14814 48242
rect 14866 48190 14868 48242
rect 14812 48132 14868 48190
rect 14812 48066 14868 48076
rect 14924 51324 15092 51380
rect 14924 47570 14980 51324
rect 15036 50708 15092 50718
rect 15036 50614 15092 50652
rect 15260 50036 15316 50046
rect 15260 49942 15316 49980
rect 15260 49588 15316 49598
rect 15260 48804 15316 49532
rect 14924 47518 14926 47570
rect 14978 47518 14980 47570
rect 14924 47506 14980 47518
rect 15148 48802 15316 48804
rect 15148 48750 15262 48802
rect 15314 48750 15316 48802
rect 15148 48748 15316 48750
rect 14588 46734 14590 46786
rect 14642 46734 14644 46786
rect 14588 46722 14644 46734
rect 15148 46564 15204 48748
rect 15260 48738 15316 48748
rect 15372 48468 15428 53678
rect 15484 53172 15540 54350
rect 15708 53732 15764 53742
rect 15708 53638 15764 53676
rect 15932 53730 15988 53742
rect 15932 53678 15934 53730
rect 15986 53678 15988 53730
rect 15484 52052 15540 53116
rect 15932 52946 15988 53678
rect 15932 52894 15934 52946
rect 15986 52894 15988 52946
rect 15484 51986 15540 51996
rect 15820 52162 15876 52174
rect 15820 52110 15822 52162
rect 15874 52110 15876 52162
rect 15484 51492 15540 51502
rect 15484 51378 15540 51436
rect 15484 51326 15486 51378
rect 15538 51326 15540 51378
rect 15484 51314 15540 51326
rect 15596 51156 15652 51166
rect 15820 51156 15876 52110
rect 15596 51154 15876 51156
rect 15596 51102 15598 51154
rect 15650 51102 15876 51154
rect 15596 51100 15876 51102
rect 15596 51090 15652 51100
rect 15932 50708 15988 52894
rect 16044 52724 16100 55918
rect 16268 54404 16324 54414
rect 16268 54310 16324 54348
rect 16380 53954 16436 57148
rect 18284 56644 18340 56654
rect 18172 56308 18228 56318
rect 17836 56196 17892 56206
rect 16492 55972 16548 55982
rect 17500 55972 17556 55982
rect 16492 55970 16772 55972
rect 16492 55918 16494 55970
rect 16546 55918 16772 55970
rect 16492 55916 16772 55918
rect 16492 55858 16548 55916
rect 16492 55806 16494 55858
rect 16546 55806 16548 55858
rect 16492 55794 16548 55806
rect 16604 55300 16660 55310
rect 16380 53902 16382 53954
rect 16434 53902 16436 53954
rect 16380 53890 16436 53902
rect 16492 55186 16548 55198
rect 16492 55134 16494 55186
rect 16546 55134 16548 55186
rect 16492 55076 16548 55134
rect 16492 53956 16548 55020
rect 16604 54514 16660 55244
rect 16716 54628 16772 55916
rect 17276 55970 17556 55972
rect 17276 55918 17502 55970
rect 17554 55918 17556 55970
rect 17276 55916 17556 55918
rect 17164 55074 17220 55086
rect 17164 55022 17166 55074
rect 17218 55022 17220 55074
rect 16716 54562 16772 54572
rect 16828 54626 16884 54638
rect 16828 54574 16830 54626
rect 16882 54574 16884 54626
rect 16604 54462 16606 54514
rect 16658 54462 16660 54514
rect 16604 54450 16660 54462
rect 16380 52836 16436 52846
rect 16380 52742 16436 52780
rect 16044 52658 16100 52668
rect 16156 52164 16212 52174
rect 16156 52070 16212 52108
rect 15596 50652 15988 50708
rect 16156 51492 16212 51502
rect 15596 50596 15652 50652
rect 15596 50502 15652 50540
rect 16044 50594 16100 50606
rect 16044 50542 16046 50594
rect 16098 50542 16100 50594
rect 15820 49700 15876 49710
rect 15820 49698 15988 49700
rect 15820 49646 15822 49698
rect 15874 49646 15988 49698
rect 15820 49644 15988 49646
rect 15820 49634 15876 49644
rect 15708 49028 15764 49038
rect 15708 48934 15764 48972
rect 15372 48402 15428 48412
rect 15820 48916 15876 48926
rect 15260 48242 15316 48254
rect 15260 48190 15262 48242
rect 15314 48190 15316 48242
rect 15260 47348 15316 48190
rect 15596 48244 15652 48254
rect 15596 48150 15652 48188
rect 15820 47460 15876 48860
rect 15820 47366 15876 47404
rect 15260 47292 15652 47348
rect 15484 47124 15540 47134
rect 15372 47068 15484 47124
rect 15260 46564 15316 46574
rect 15148 46508 15260 46564
rect 14252 46450 14420 46452
rect 14252 46398 14254 46450
rect 14306 46398 14420 46450
rect 14252 46396 14420 46398
rect 14812 46450 14868 46462
rect 15036 46452 15092 46462
rect 14812 46398 14814 46450
rect 14866 46398 14868 46450
rect 14140 45890 14196 45902
rect 14140 45838 14142 45890
rect 14194 45838 14196 45890
rect 14140 45780 14196 45838
rect 14252 45892 14308 46396
rect 14364 45892 14420 45902
rect 14252 45890 14420 45892
rect 14252 45838 14366 45890
rect 14418 45838 14420 45890
rect 14252 45836 14420 45838
rect 14364 45826 14420 45836
rect 14140 45714 14196 45724
rect 14140 45444 14196 45454
rect 14028 45218 14084 45230
rect 14028 45166 14030 45218
rect 14082 45166 14084 45218
rect 14028 44324 14084 45166
rect 14140 44994 14196 45388
rect 14812 45444 14868 46398
rect 14812 45378 14868 45388
rect 14924 46450 15092 46452
rect 14924 46398 15038 46450
rect 15090 46398 15092 46450
rect 14924 46396 15092 46398
rect 14140 44942 14142 44994
rect 14194 44942 14196 44994
rect 14140 44930 14196 44942
rect 14924 44994 14980 46396
rect 15036 46386 15092 46396
rect 14924 44942 14926 44994
rect 14978 44942 14980 44994
rect 14812 44548 14868 44558
rect 14812 44454 14868 44492
rect 14924 44324 14980 44942
rect 14084 44268 14196 44324
rect 14028 44258 14084 44268
rect 14028 44100 14084 44110
rect 14028 44006 14084 44044
rect 13916 43820 14084 43876
rect 13916 43538 13972 43550
rect 13916 43486 13918 43538
rect 13970 43486 13972 43538
rect 13804 42756 13860 42766
rect 13356 41794 13412 41804
rect 13468 42754 13860 42756
rect 13468 42702 13806 42754
rect 13858 42702 13860 42754
rect 13468 42700 13860 42702
rect 13468 42082 13524 42700
rect 13804 42690 13860 42700
rect 13916 42420 13972 43486
rect 13468 42030 13470 42082
rect 13522 42030 13524 42082
rect 13468 41186 13524 42030
rect 13468 41134 13470 41186
rect 13522 41134 13524 41186
rect 13468 41122 13524 41134
rect 13804 42364 13972 42420
rect 13804 41972 13860 42364
rect 13916 42196 13972 42206
rect 14028 42196 14084 43820
rect 14140 43540 14196 44268
rect 14588 44268 14980 44324
rect 15260 44994 15316 46508
rect 15260 44942 15262 44994
rect 15314 44942 15316 44994
rect 14476 44210 14532 44222
rect 14476 44158 14478 44210
rect 14530 44158 14532 44210
rect 14476 44100 14532 44158
rect 14476 44034 14532 44044
rect 14364 43652 14420 43662
rect 14364 43558 14420 43596
rect 14140 43474 14196 43484
rect 14588 43428 14644 44268
rect 14700 44100 14756 44110
rect 14700 43764 14756 44044
rect 15148 44100 15204 44110
rect 15148 44006 15204 44044
rect 14700 43698 14756 43708
rect 14924 43650 14980 43662
rect 14924 43598 14926 43650
rect 14978 43598 14980 43650
rect 13916 42194 14084 42196
rect 13916 42142 13918 42194
rect 13970 42142 14084 42194
rect 13916 42140 14084 42142
rect 14252 43372 14644 43428
rect 14812 43538 14868 43550
rect 14812 43486 14814 43538
rect 14866 43486 14868 43538
rect 13916 42130 13972 42140
rect 13692 40404 13748 40414
rect 13804 40404 13860 41916
rect 14252 41074 14308 43372
rect 14588 41972 14644 41982
rect 14812 41972 14868 43486
rect 14924 43540 14980 43598
rect 14980 43484 15204 43540
rect 14924 43474 14980 43484
rect 14924 43314 14980 43326
rect 14924 43262 14926 43314
rect 14978 43262 14980 43314
rect 14924 42196 14980 43262
rect 14924 42130 14980 42140
rect 15036 42754 15092 42766
rect 15036 42702 15038 42754
rect 15090 42702 15092 42754
rect 14924 41972 14980 41982
rect 14812 41916 14924 41972
rect 14588 41878 14644 41916
rect 14924 41878 14980 41916
rect 14364 41188 14420 41198
rect 14812 41188 14868 41198
rect 15036 41188 15092 42702
rect 15148 42084 15204 43484
rect 15260 42308 15316 44942
rect 15372 43204 15428 47068
rect 15484 47058 15540 47068
rect 15484 46004 15540 46014
rect 15484 45890 15540 45948
rect 15484 45838 15486 45890
rect 15538 45838 15540 45890
rect 15484 44436 15540 45838
rect 15484 44370 15540 44380
rect 15596 45890 15652 47292
rect 15932 46340 15988 49644
rect 16044 47908 16100 50542
rect 16044 47842 16100 47852
rect 16156 47684 16212 51436
rect 16380 51378 16436 51390
rect 16380 51326 16382 51378
rect 16434 51326 16436 51378
rect 16380 51268 16436 51326
rect 16380 50484 16436 51212
rect 16380 50418 16436 50428
rect 16268 49700 16324 49710
rect 16268 49026 16324 49644
rect 16268 48974 16270 49026
rect 16322 48974 16324 49026
rect 16268 48962 16324 48974
rect 16380 49698 16436 49710
rect 16380 49646 16382 49698
rect 16434 49646 16436 49698
rect 16380 48916 16436 49646
rect 16380 48850 16436 48860
rect 16156 47618 16212 47628
rect 16380 47460 16436 47470
rect 16156 47458 16436 47460
rect 16156 47406 16382 47458
rect 16434 47406 16436 47458
rect 16156 47404 16436 47406
rect 16044 47012 16100 47022
rect 16044 46898 16100 46956
rect 16044 46846 16046 46898
rect 16098 46846 16100 46898
rect 16044 46834 16100 46846
rect 15932 46274 15988 46284
rect 15596 45838 15598 45890
rect 15650 45838 15652 45890
rect 15484 43988 15540 43998
rect 15484 43316 15540 43932
rect 15596 43540 15652 45838
rect 15708 46114 15764 46126
rect 15708 46062 15710 46114
rect 15762 46062 15764 46114
rect 15708 45892 15764 46062
rect 15932 45892 15988 45902
rect 15708 45890 15988 45892
rect 15708 45838 15934 45890
rect 15986 45838 15988 45890
rect 15708 45836 15988 45838
rect 15932 45826 15988 45836
rect 15708 44994 15764 45006
rect 15708 44942 15710 44994
rect 15762 44942 15764 44994
rect 15708 44884 15764 44942
rect 15708 44818 15764 44828
rect 15820 44660 15876 44670
rect 15708 44324 15764 44334
rect 15708 44230 15764 44268
rect 15596 43474 15652 43484
rect 15708 43426 15764 43438
rect 15708 43374 15710 43426
rect 15762 43374 15764 43426
rect 15708 43316 15764 43374
rect 15484 43260 15764 43316
rect 15372 43148 15652 43204
rect 15260 42242 15316 42252
rect 15484 42084 15540 42094
rect 15148 42082 15540 42084
rect 15148 42030 15486 42082
rect 15538 42030 15540 42082
rect 15148 42028 15540 42030
rect 15484 42018 15540 42028
rect 14364 41094 14420 41132
rect 14588 41186 15092 41188
rect 14588 41134 14814 41186
rect 14866 41134 15092 41186
rect 14588 41132 15092 41134
rect 15148 41860 15204 41870
rect 14252 41022 14254 41074
rect 14306 41022 14308 41074
rect 13692 40402 13860 40404
rect 13692 40350 13694 40402
rect 13746 40350 13860 40402
rect 13692 40348 13860 40350
rect 14140 40404 14196 40414
rect 13468 39732 13524 39742
rect 12908 39564 13076 39620
rect 13020 38668 13076 39564
rect 13468 39618 13524 39676
rect 13468 39566 13470 39618
rect 13522 39566 13524 39618
rect 13468 39058 13524 39566
rect 13468 39006 13470 39058
rect 13522 39006 13524 39058
rect 13468 38994 13524 39006
rect 12684 37102 12686 37154
rect 12738 37102 12740 37154
rect 12684 37090 12740 37102
rect 12908 38612 13076 38668
rect 13132 38724 13188 38734
rect 13132 38630 13188 38668
rect 11788 36502 11844 36540
rect 12124 36482 12180 36494
rect 12124 36430 12126 36482
rect 12178 36430 12180 36482
rect 12124 36260 12180 36430
rect 12348 36484 12404 36494
rect 12348 36390 12404 36428
rect 11116 36082 11172 36092
rect 11900 36204 12180 36260
rect 12908 36370 12964 38612
rect 13468 37828 13524 37838
rect 13468 37734 13524 37772
rect 13692 37380 13748 40348
rect 14028 39618 14084 39630
rect 14028 39566 14030 39618
rect 14082 39566 14084 39618
rect 14028 39508 14084 39566
rect 14028 39442 14084 39452
rect 14028 38836 14084 38846
rect 14140 38836 14196 40348
rect 14028 38834 14196 38836
rect 14028 38782 14030 38834
rect 14082 38782 14196 38834
rect 14028 38780 14196 38782
rect 14028 38770 14084 38780
rect 14252 38388 14308 41022
rect 14588 39506 14644 41132
rect 14812 41122 14868 41132
rect 14924 40628 14980 40638
rect 15148 40628 15204 41804
rect 14980 40572 15092 40628
rect 14924 40562 14980 40572
rect 14700 40404 14756 40414
rect 14700 39618 14756 40348
rect 14812 40402 14868 40414
rect 14812 40350 14814 40402
rect 14866 40350 14868 40402
rect 14812 40180 14868 40350
rect 14812 40114 14868 40124
rect 14924 40178 14980 40190
rect 14924 40126 14926 40178
rect 14978 40126 14980 40178
rect 14924 39956 14980 40126
rect 14924 39890 14980 39900
rect 14700 39566 14702 39618
rect 14754 39566 14756 39618
rect 14700 39554 14756 39566
rect 14924 39732 14980 39742
rect 14588 39454 14590 39506
rect 14642 39454 14644 39506
rect 14588 39060 14644 39454
rect 14812 39508 14868 39518
rect 14476 39004 14644 39060
rect 14700 39284 14756 39294
rect 14364 38948 14420 38958
rect 14364 38668 14420 38892
rect 14476 38668 14532 39004
rect 14700 38668 14756 39228
rect 14812 38834 14868 39452
rect 14924 39172 14980 39676
rect 14924 39106 14980 39116
rect 14812 38782 14814 38834
rect 14866 38782 14868 38834
rect 14812 38770 14868 38782
rect 15036 38668 15092 40572
rect 15148 40562 15204 40572
rect 15372 41300 15428 41310
rect 15372 39618 15428 41244
rect 15372 39566 15374 39618
rect 15426 39566 15428 39618
rect 15372 39554 15428 39566
rect 15484 39396 15540 39406
rect 15596 39396 15652 43148
rect 15708 42756 15764 43260
rect 15708 42690 15764 42700
rect 15820 42532 15876 44604
rect 16156 43538 16212 47404
rect 16380 47394 16436 47404
rect 16380 47236 16436 47246
rect 16268 46788 16324 46826
rect 16268 46722 16324 46732
rect 16380 46002 16436 47180
rect 16492 46900 16548 53900
rect 16716 51268 16772 51278
rect 16604 51266 16772 51268
rect 16604 51214 16718 51266
rect 16770 51214 16772 51266
rect 16604 51212 16772 51214
rect 16604 50428 16660 51212
rect 16716 51202 16772 51212
rect 16828 51156 16884 54574
rect 17052 54292 17108 54302
rect 17052 54068 17108 54236
rect 17052 54002 17108 54012
rect 16940 53732 16996 53742
rect 16940 53730 17108 53732
rect 16940 53678 16942 53730
rect 16994 53678 17108 53730
rect 16940 53676 17108 53678
rect 16940 53666 16996 53676
rect 16828 51090 16884 51100
rect 17052 52500 17108 53676
rect 17164 53508 17220 55022
rect 17164 53442 17220 53452
rect 17276 52836 17332 55916
rect 17500 55906 17556 55916
rect 17836 55972 17892 56140
rect 17836 55410 17892 55916
rect 17836 55358 17838 55410
rect 17890 55358 17892 55410
rect 17836 55346 17892 55358
rect 17948 55970 18004 55982
rect 17948 55918 17950 55970
rect 18002 55918 18004 55970
rect 17388 55188 17444 55198
rect 17388 54068 17444 55132
rect 17500 55074 17556 55086
rect 17500 55022 17502 55074
rect 17554 55022 17556 55074
rect 17500 54516 17556 55022
rect 17724 54516 17780 54526
rect 17500 54514 17780 54516
rect 17500 54462 17726 54514
rect 17778 54462 17780 54514
rect 17500 54460 17780 54462
rect 17724 54450 17780 54460
rect 17836 54516 17892 54526
rect 17388 54002 17444 54012
rect 17276 52770 17332 52780
rect 17388 53618 17444 53630
rect 17388 53566 17390 53618
rect 17442 53566 17444 53618
rect 16716 50932 16772 50942
rect 16716 50706 16772 50876
rect 16716 50654 16718 50706
rect 16770 50654 16772 50706
rect 16716 50642 16772 50654
rect 16940 50820 16996 50830
rect 16940 50594 16996 50764
rect 16940 50542 16942 50594
rect 16994 50542 16996 50594
rect 16940 50530 16996 50542
rect 17052 50428 17108 52444
rect 17164 52612 17220 52622
rect 17164 52050 17220 52556
rect 17164 51998 17166 52050
rect 17218 51998 17220 52050
rect 17164 51986 17220 51998
rect 16604 50372 16772 50428
rect 17052 50372 17332 50428
rect 16604 50148 16660 50158
rect 16604 48804 16660 50092
rect 16604 47124 16660 48748
rect 16716 48692 16772 50372
rect 16828 50260 16884 50270
rect 16828 50034 16884 50204
rect 16828 49982 16830 50034
rect 16882 49982 16884 50034
rect 16828 49924 16884 49982
rect 16828 49858 16884 49868
rect 16828 49138 16884 49150
rect 16828 49086 16830 49138
rect 16882 49086 16884 49138
rect 16828 49028 16884 49086
rect 16828 48962 16884 48972
rect 16940 49026 16996 49038
rect 16940 48974 16942 49026
rect 16994 48974 16996 49026
rect 16716 48626 16772 48636
rect 16828 48356 16884 48366
rect 16828 47460 16884 48300
rect 16716 47348 16772 47358
rect 16828 47348 16884 47404
rect 16716 47346 16884 47348
rect 16716 47294 16718 47346
rect 16770 47294 16884 47346
rect 16716 47292 16884 47294
rect 16716 47282 16772 47292
rect 16604 47068 16772 47124
rect 16492 46834 16548 46844
rect 16492 46564 16548 46574
rect 16492 46470 16548 46508
rect 16716 46228 16772 47068
rect 16828 46900 16884 46910
rect 16828 46806 16884 46844
rect 16380 45950 16382 46002
rect 16434 45950 16436 46002
rect 16380 45938 16436 45950
rect 16492 46172 16772 46228
rect 16828 46228 16884 46238
rect 16380 44994 16436 45006
rect 16380 44942 16382 44994
rect 16434 44942 16436 44994
rect 16380 44324 16436 44942
rect 16380 44258 16436 44268
rect 16156 43486 16158 43538
rect 16210 43486 16212 43538
rect 15372 39394 15652 39396
rect 15372 39342 15486 39394
rect 15538 39342 15652 39394
rect 15372 39340 15652 39342
rect 15708 42476 15876 42532
rect 16044 42754 16100 42766
rect 16044 42702 16046 42754
rect 16098 42702 16100 42754
rect 15260 39060 15316 39070
rect 15260 38834 15316 39004
rect 15260 38782 15262 38834
rect 15314 38782 15316 38834
rect 15260 38770 15316 38782
rect 14364 38612 14532 38668
rect 14252 38322 14308 38332
rect 14476 38164 14532 38612
rect 14588 38612 14756 38668
rect 14812 38612 15092 38668
rect 15372 38612 15428 39340
rect 15484 39330 15540 39340
rect 15708 39284 15764 42476
rect 16044 41186 16100 42702
rect 16156 42644 16212 43486
rect 16156 42578 16212 42588
rect 16268 44212 16324 44222
rect 16268 42642 16324 44156
rect 16268 42590 16270 42642
rect 16322 42590 16324 42642
rect 16268 41524 16324 42590
rect 16268 41458 16324 41468
rect 16380 43428 16436 43438
rect 16044 41134 16046 41186
rect 16098 41134 16100 41186
rect 15820 40404 15876 40414
rect 16044 40404 16100 41134
rect 15820 40402 16100 40404
rect 15820 40350 15822 40402
rect 15874 40350 16100 40402
rect 15820 40348 16100 40350
rect 16268 41188 16324 41198
rect 16268 40626 16324 41132
rect 16268 40574 16270 40626
rect 16322 40574 16324 40626
rect 16268 40404 16324 40574
rect 16380 40626 16436 43372
rect 16492 43426 16548 46172
rect 16828 45892 16884 46172
rect 16492 43374 16494 43426
rect 16546 43374 16548 43426
rect 16492 43362 16548 43374
rect 16604 45836 16884 45892
rect 16604 44322 16660 45836
rect 16716 45220 16772 45230
rect 16716 44548 16772 45164
rect 16716 44434 16772 44492
rect 16716 44382 16718 44434
rect 16770 44382 16772 44434
rect 16716 44370 16772 44382
rect 16828 44994 16884 45006
rect 16828 44942 16830 44994
rect 16882 44942 16884 44994
rect 16828 44884 16884 44942
rect 16604 44270 16606 44322
rect 16658 44270 16660 44322
rect 16604 42978 16660 44270
rect 16828 44212 16884 44828
rect 16940 44434 16996 48974
rect 17276 48356 17332 50372
rect 17388 50036 17444 53566
rect 17836 53618 17892 54460
rect 17836 53566 17838 53618
rect 17890 53566 17892 53618
rect 17836 53554 17892 53566
rect 17948 53508 18004 55918
rect 18060 55524 18116 55534
rect 18060 55430 18116 55468
rect 18172 54292 18228 56252
rect 18284 56306 18340 56588
rect 18284 56254 18286 56306
rect 18338 56254 18340 56306
rect 18284 56242 18340 56254
rect 19628 56644 19684 56654
rect 19180 56196 19236 56206
rect 19236 56140 19348 56196
rect 19180 56102 19236 56140
rect 19068 56082 19124 56094
rect 19068 56030 19070 56082
rect 19122 56030 19124 56082
rect 18844 55972 18900 56010
rect 18844 55906 18900 55916
rect 18844 55748 18900 55758
rect 18732 55300 18788 55310
rect 18732 55206 18788 55244
rect 18396 55074 18452 55086
rect 18396 55022 18398 55074
rect 18450 55022 18452 55074
rect 18396 54516 18452 55022
rect 18844 54516 18900 55692
rect 19068 55524 19124 56030
rect 19180 55860 19236 55870
rect 19180 55766 19236 55804
rect 19068 55458 19124 55468
rect 19180 55636 19236 55646
rect 19068 55300 19124 55310
rect 19180 55300 19236 55580
rect 19068 55298 19236 55300
rect 19068 55246 19070 55298
rect 19122 55246 19236 55298
rect 19068 55244 19236 55246
rect 19068 55234 19124 55244
rect 19068 54516 19124 54526
rect 18844 54514 19124 54516
rect 18844 54462 19070 54514
rect 19122 54462 19124 54514
rect 18844 54460 19124 54462
rect 18396 54450 18452 54460
rect 19068 54450 19124 54460
rect 18172 53954 18228 54236
rect 18172 53902 18174 53954
rect 18226 53902 18228 53954
rect 18172 53890 18228 53902
rect 18060 53844 18116 53854
rect 18060 53750 18116 53788
rect 18844 53508 18900 53518
rect 17948 53452 18228 53508
rect 17500 53396 17556 53406
rect 17500 53172 17556 53340
rect 17500 53078 17556 53116
rect 17836 53284 17892 53294
rect 17612 52276 17668 52286
rect 17612 52182 17668 52220
rect 17724 51380 17780 51390
rect 17500 50596 17556 50606
rect 17500 50502 17556 50540
rect 17724 50428 17780 51324
rect 17836 51380 17892 53228
rect 18060 52834 18116 52846
rect 18060 52782 18062 52834
rect 18114 52782 18116 52834
rect 18060 52388 18116 52782
rect 18060 52322 18116 52332
rect 18060 51940 18116 51950
rect 18172 51940 18228 53452
rect 18844 53170 18900 53452
rect 18844 53118 18846 53170
rect 18898 53118 18900 53170
rect 18844 53106 18900 53118
rect 18508 52948 18564 52958
rect 18508 52946 18788 52948
rect 18508 52894 18510 52946
rect 18562 52894 18788 52946
rect 18508 52892 18788 52894
rect 18508 52882 18564 52892
rect 18620 52724 18676 52734
rect 18284 52612 18340 52622
rect 18284 52274 18340 52556
rect 18284 52222 18286 52274
rect 18338 52222 18340 52274
rect 18284 52052 18340 52222
rect 18620 52164 18676 52668
rect 18284 51986 18340 51996
rect 18396 52162 18676 52164
rect 18396 52110 18622 52162
rect 18674 52110 18676 52162
rect 18396 52108 18676 52110
rect 18116 51884 18228 51940
rect 18060 51874 18116 51884
rect 18060 51492 18116 51502
rect 17948 51380 18004 51390
rect 17836 51324 17948 51380
rect 17836 51266 17892 51324
rect 17948 51314 18004 51324
rect 17836 51214 17838 51266
rect 17890 51214 17892 51266
rect 17836 51202 17892 51214
rect 18060 50596 18116 51436
rect 18396 50820 18452 52108
rect 18620 52098 18676 52108
rect 18732 51604 18788 52892
rect 19180 52946 19236 52958
rect 19180 52894 19182 52946
rect 19234 52894 19236 52946
rect 19180 52276 19236 52894
rect 19180 52210 19236 52220
rect 19292 51716 19348 56140
rect 19628 55410 19684 56588
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 21084 56306 21140 57260
rect 21084 56254 21086 56306
rect 21138 56254 21140 56306
rect 21084 56242 21140 56254
rect 20972 56196 21028 56206
rect 19740 56082 19796 56094
rect 19740 56030 19742 56082
rect 19794 56030 19796 56082
rect 19740 55524 19796 56030
rect 20188 56084 20244 56094
rect 20412 56084 20468 56094
rect 19740 55458 19796 55468
rect 20076 55970 20132 55982
rect 20076 55918 20078 55970
rect 20130 55918 20132 55970
rect 19628 55358 19630 55410
rect 19682 55358 19684 55410
rect 19628 54292 19684 55358
rect 20076 55076 20132 55918
rect 20188 55300 20244 56028
rect 20188 55234 20244 55244
rect 20300 56028 20412 56084
rect 20076 55020 20244 55076
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 20188 54740 20244 55020
rect 20076 54684 20244 54740
rect 19740 54516 19796 54526
rect 19740 54422 19796 54460
rect 19628 54236 19796 54292
rect 19628 54068 19684 54078
rect 19404 53956 19460 53966
rect 19404 53862 19460 53900
rect 19628 53730 19684 54012
rect 19628 53678 19630 53730
rect 19682 53678 19684 53730
rect 19628 53666 19684 53678
rect 19740 53508 19796 54236
rect 19628 53452 19796 53508
rect 20076 53508 20132 54684
rect 20076 53452 20244 53508
rect 19404 53060 19460 53070
rect 19404 52386 19460 53004
rect 19404 52334 19406 52386
rect 19458 52334 19460 52386
rect 19404 52322 19460 52334
rect 19628 52276 19684 53452
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 19740 52946 19796 52958
rect 19740 52894 19742 52946
rect 19794 52894 19796 52946
rect 19740 52836 19796 52894
rect 19740 52770 19796 52780
rect 20188 52836 20244 53452
rect 20188 52770 20244 52780
rect 20300 52388 20356 56028
rect 20412 56018 20468 56028
rect 20748 55412 20804 55422
rect 20748 55300 20804 55356
rect 20524 55298 20804 55300
rect 20524 55246 20750 55298
rect 20802 55246 20804 55298
rect 20524 55244 20804 55246
rect 20412 53844 20468 53854
rect 20412 53750 20468 53788
rect 20524 53730 20580 55244
rect 20748 55234 20804 55244
rect 20524 53678 20526 53730
rect 20578 53678 20580 53730
rect 20524 53666 20580 53678
rect 20860 54626 20916 54638
rect 20860 54574 20862 54626
rect 20914 54574 20916 54626
rect 20636 53508 20692 53518
rect 19628 52210 19684 52220
rect 20188 52332 20356 52388
rect 20524 53506 20692 53508
rect 20524 53454 20638 53506
rect 20690 53454 20692 53506
rect 20524 53452 20692 53454
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19292 51660 19684 51716
rect 19836 51706 20100 51716
rect 19628 51604 19684 51660
rect 19628 51548 19796 51604
rect 18732 51538 18788 51548
rect 18844 51378 18900 51390
rect 18844 51326 18846 51378
rect 18898 51326 18900 51378
rect 18844 51268 18900 51326
rect 19180 51380 19236 51390
rect 19180 51286 19236 51324
rect 19628 51378 19684 51390
rect 19628 51326 19630 51378
rect 19682 51326 19684 51378
rect 17388 49970 17444 49980
rect 17612 50372 17780 50428
rect 17836 50482 17892 50494
rect 18060 50484 18116 50540
rect 17836 50430 17838 50482
rect 17890 50430 17892 50482
rect 17276 48290 17332 48300
rect 17388 49812 17444 49822
rect 17388 48132 17444 49756
rect 17500 49028 17556 49038
rect 17500 48934 17556 48972
rect 17276 48076 17444 48132
rect 17052 47572 17108 47582
rect 17052 47478 17108 47516
rect 17276 47460 17332 48076
rect 17164 47458 17332 47460
rect 17164 47406 17278 47458
rect 17330 47406 17332 47458
rect 17164 47404 17332 47406
rect 16940 44382 16942 44434
rect 16994 44382 16996 44434
rect 16940 44370 16996 44382
rect 17052 46676 17108 46686
rect 16828 44146 16884 44156
rect 16604 42926 16606 42978
rect 16658 42926 16660 42978
rect 16604 42914 16660 42926
rect 17052 42868 17108 46620
rect 16940 42812 17108 42868
rect 16940 40740 16996 42812
rect 16940 40674 16996 40684
rect 17052 42644 17108 42654
rect 17164 42644 17220 47404
rect 17276 47394 17332 47404
rect 17388 47460 17444 47470
rect 17388 46674 17444 47404
rect 17388 46622 17390 46674
rect 17442 46622 17444 46674
rect 17388 46610 17444 46622
rect 17612 46676 17668 50372
rect 17724 48916 17780 48954
rect 17724 48850 17780 48860
rect 17612 46610 17668 46620
rect 17724 48692 17780 48702
rect 17724 47460 17780 48636
rect 17612 46452 17668 46462
rect 17388 46450 17668 46452
rect 17388 46398 17614 46450
rect 17666 46398 17668 46450
rect 17388 46396 17668 46398
rect 17276 44322 17332 44334
rect 17276 44270 17278 44322
rect 17330 44270 17332 44322
rect 17276 44212 17332 44270
rect 17276 44146 17332 44156
rect 17388 43652 17444 46396
rect 17612 46386 17668 46396
rect 17612 46114 17668 46126
rect 17612 46062 17614 46114
rect 17666 46062 17668 46114
rect 17500 46002 17556 46014
rect 17500 45950 17502 46002
rect 17554 45950 17556 46002
rect 17500 45556 17556 45950
rect 17500 45490 17556 45500
rect 17500 45330 17556 45342
rect 17500 45278 17502 45330
rect 17554 45278 17556 45330
rect 17500 45108 17556 45278
rect 17612 45330 17668 46062
rect 17612 45278 17614 45330
rect 17666 45278 17668 45330
rect 17612 45266 17668 45278
rect 17724 45108 17780 47404
rect 17836 46228 17892 50430
rect 17948 50428 18116 50484
rect 18284 50764 18452 50820
rect 18620 51154 18676 51166
rect 18620 51102 18622 51154
rect 18674 51102 18676 51154
rect 18284 50428 18340 50764
rect 18396 50596 18452 50606
rect 18620 50596 18676 51102
rect 18396 50594 18620 50596
rect 18396 50542 18398 50594
rect 18450 50542 18620 50594
rect 18396 50540 18620 50542
rect 18396 50530 18452 50540
rect 18620 50530 18676 50540
rect 18732 51156 18788 51166
rect 18732 50708 18788 51100
rect 18732 50594 18788 50652
rect 18732 50542 18734 50594
rect 18786 50542 18788 50594
rect 18732 50530 18788 50542
rect 17948 49810 18004 50428
rect 18284 50372 18452 50428
rect 17948 49758 17950 49810
rect 18002 49758 18004 49810
rect 17948 49746 18004 49758
rect 18284 49700 18340 49710
rect 18284 49606 18340 49644
rect 17948 47908 18004 47918
rect 17948 46674 18004 47852
rect 18284 47796 18340 47806
rect 18172 47740 18284 47796
rect 18060 47458 18116 47470
rect 18060 47406 18062 47458
rect 18114 47406 18116 47458
rect 18060 47124 18116 47406
rect 18060 47058 18116 47068
rect 18172 47012 18228 47740
rect 18284 47730 18340 47740
rect 18284 47458 18340 47470
rect 18284 47406 18286 47458
rect 18338 47406 18340 47458
rect 18284 47348 18340 47406
rect 18284 47282 18340 47292
rect 17948 46622 17950 46674
rect 18002 46622 18004 46674
rect 17948 46610 18004 46622
rect 18060 46900 18116 46910
rect 18172 46900 18228 46956
rect 18060 46898 18228 46900
rect 18060 46846 18062 46898
rect 18114 46846 18228 46898
rect 18060 46844 18228 46846
rect 17836 46162 17892 46172
rect 17500 45052 17780 45108
rect 17836 45778 17892 45790
rect 17836 45726 17838 45778
rect 17890 45726 17892 45778
rect 17724 44882 17780 44894
rect 17724 44830 17726 44882
rect 17778 44830 17780 44882
rect 17724 44660 17780 44830
rect 17724 44594 17780 44604
rect 17612 44212 17668 44222
rect 17108 42588 17220 42644
rect 17276 43596 17444 43652
rect 17500 44210 17668 44212
rect 17500 44158 17614 44210
rect 17666 44158 17668 44210
rect 17500 44156 17668 44158
rect 16380 40574 16382 40626
rect 16434 40574 16436 40626
rect 16380 40562 16436 40574
rect 16492 40628 16548 40638
rect 16492 40534 16548 40572
rect 15820 40292 15876 40348
rect 16268 40338 16324 40348
rect 16940 40402 16996 40414
rect 16940 40350 16942 40402
rect 16994 40350 16996 40402
rect 16940 40292 16996 40350
rect 15820 39620 15876 40236
rect 16828 40236 16940 40292
rect 15820 39554 15876 39564
rect 16268 39732 16324 39742
rect 15596 39228 15764 39284
rect 15596 38668 15652 39228
rect 14588 38610 14644 38612
rect 14588 38558 14590 38610
rect 14642 38558 14644 38610
rect 14588 38546 14644 38558
rect 14812 38276 14868 38612
rect 15372 38546 15428 38556
rect 15484 38612 15652 38668
rect 16268 39058 16324 39676
rect 16604 39620 16660 39630
rect 16604 39526 16660 39564
rect 16268 39006 16270 39058
rect 16322 39006 16324 39058
rect 15484 38388 15540 38612
rect 14700 38274 14868 38276
rect 14700 38222 14814 38274
rect 14866 38222 14868 38274
rect 14700 38220 14868 38222
rect 14588 38164 14644 38174
rect 14476 38162 14644 38164
rect 14476 38110 14590 38162
rect 14642 38110 14644 38162
rect 14476 38108 14644 38110
rect 14588 38098 14644 38108
rect 14028 38050 14084 38062
rect 14028 37998 14030 38050
rect 14082 37998 14084 38050
rect 14028 37940 14084 37998
rect 14700 37940 14756 38220
rect 14812 38210 14868 38220
rect 15148 38332 15540 38388
rect 15148 38274 15204 38332
rect 15148 38222 15150 38274
rect 15202 38222 15204 38274
rect 15148 38210 15204 38222
rect 16156 38164 16212 38174
rect 16156 38070 16212 38108
rect 16268 38052 16324 39006
rect 16828 38946 16884 40236
rect 16940 40226 16996 40236
rect 16940 39618 16996 39630
rect 16940 39566 16942 39618
rect 16994 39566 16996 39618
rect 16940 39508 16996 39566
rect 16940 39442 16996 39452
rect 16828 38894 16830 38946
rect 16882 38894 16884 38946
rect 16828 38882 16884 38894
rect 17052 38162 17108 42588
rect 17164 42420 17220 42430
rect 17164 41410 17220 42364
rect 17164 41358 17166 41410
rect 17218 41358 17220 41410
rect 17164 41346 17220 41358
rect 17052 38110 17054 38162
rect 17106 38110 17108 38162
rect 17052 38098 17108 38110
rect 17164 41186 17220 41198
rect 17164 41134 17166 41186
rect 17218 41134 17220 41186
rect 17164 38836 17220 41134
rect 17276 41076 17332 43596
rect 17388 43428 17444 43438
rect 17388 43334 17444 43372
rect 17388 41972 17444 41982
rect 17388 41878 17444 41916
rect 17500 41860 17556 44156
rect 17612 44146 17668 44156
rect 17724 44212 17780 44222
rect 17500 41794 17556 41804
rect 17612 43988 17668 43998
rect 17612 42754 17668 43932
rect 17724 43764 17780 44156
rect 17724 43538 17780 43708
rect 17724 43486 17726 43538
rect 17778 43486 17780 43538
rect 17724 43474 17780 43486
rect 17612 42702 17614 42754
rect 17666 42702 17668 42754
rect 17388 41412 17444 41422
rect 17388 41188 17444 41356
rect 17388 41094 17444 41132
rect 17276 41010 17332 41020
rect 17276 40740 17332 40750
rect 17332 40684 17444 40740
rect 17276 40674 17332 40684
rect 17388 40290 17444 40684
rect 17388 40238 17390 40290
rect 17442 40238 17444 40290
rect 17388 40180 17444 40238
rect 17388 40114 17444 40124
rect 17164 38164 17220 38780
rect 17612 38668 17668 42702
rect 17836 41636 17892 45726
rect 18060 45444 18116 46844
rect 18172 46676 18228 46686
rect 18172 46582 18228 46620
rect 18284 46674 18340 46686
rect 18284 46622 18286 46674
rect 18338 46622 18340 46674
rect 18060 45378 18116 45388
rect 18284 45220 18340 46622
rect 18284 45154 18340 45164
rect 18284 44996 18340 45006
rect 18060 44994 18340 44996
rect 18060 44942 18286 44994
rect 18338 44942 18340 44994
rect 18060 44940 18340 44942
rect 18060 43988 18116 44940
rect 18284 44930 18340 44940
rect 18060 43922 18116 43932
rect 18396 43876 18452 50372
rect 18732 50372 18788 50382
rect 18732 50278 18788 50316
rect 18844 50148 18900 51212
rect 19628 50932 19684 51326
rect 18844 50082 18900 50092
rect 19516 50876 19684 50932
rect 18732 50036 18788 50046
rect 18732 49922 18788 49980
rect 18732 49870 18734 49922
rect 18786 49870 18788 49922
rect 18732 49858 18788 49870
rect 18508 49810 18564 49822
rect 18508 49758 18510 49810
rect 18562 49758 18564 49810
rect 18508 48804 18564 49758
rect 19292 49812 19348 49822
rect 19292 49718 19348 49756
rect 19180 49364 19236 49374
rect 19180 49026 19236 49308
rect 19180 48974 19182 49026
rect 19234 48974 19236 49026
rect 19180 48962 19236 48974
rect 18508 48738 18564 48748
rect 18732 48916 18788 48926
rect 18620 48242 18676 48254
rect 18620 48190 18622 48242
rect 18674 48190 18676 48242
rect 18508 48130 18564 48142
rect 18508 48078 18510 48130
rect 18562 48078 18564 48130
rect 18508 46900 18564 48078
rect 18620 47572 18676 48190
rect 18732 48244 18788 48860
rect 19516 48468 19572 50876
rect 19628 50596 19684 50606
rect 19628 50502 19684 50540
rect 19740 50482 19796 51548
rect 20076 51380 20132 51390
rect 20188 51380 20244 52332
rect 20300 52164 20356 52174
rect 20300 52070 20356 52108
rect 20412 52162 20468 52174
rect 20412 52110 20414 52162
rect 20466 52110 20468 52162
rect 20076 51378 20188 51380
rect 20076 51326 20078 51378
rect 20130 51326 20188 51378
rect 20076 51324 20188 51326
rect 20076 51314 20132 51324
rect 20188 51286 20244 51324
rect 20412 51268 20468 52110
rect 20412 51202 20468 51212
rect 20076 51156 20132 51166
rect 20076 51062 20132 51100
rect 20524 50932 20580 53452
rect 20636 53442 20692 53452
rect 20748 52500 20804 52510
rect 20748 52162 20804 52444
rect 20748 52110 20750 52162
rect 20802 52110 20804 52162
rect 20748 52098 20804 52110
rect 20636 51940 20692 51950
rect 20636 51846 20692 51884
rect 20860 51940 20916 54574
rect 20860 51874 20916 51884
rect 20300 50876 20580 50932
rect 20300 50594 20356 50876
rect 20300 50542 20302 50594
rect 20354 50542 20356 50594
rect 20300 50530 20356 50542
rect 19740 50430 19742 50482
rect 19794 50430 19796 50482
rect 19740 50418 19796 50430
rect 20524 50428 20580 50876
rect 20636 51492 20692 51502
rect 20636 51378 20692 51436
rect 20636 51326 20638 51378
rect 20690 51326 20692 51378
rect 20636 50932 20692 51326
rect 20748 51380 20804 51390
rect 20748 51286 20804 51324
rect 20860 51378 20916 51390
rect 20860 51326 20862 51378
rect 20914 51326 20916 51378
rect 20636 50866 20692 50876
rect 20748 50484 20804 50522
rect 19404 48412 19572 48468
rect 19628 50372 19684 50382
rect 18732 48178 18788 48188
rect 19292 48242 19348 48254
rect 19292 48190 19294 48242
rect 19346 48190 19348 48242
rect 18620 47506 18676 47516
rect 18732 48020 18788 48030
rect 18732 47012 18788 47964
rect 19180 47684 19236 47694
rect 19292 47684 19348 48190
rect 19180 47682 19348 47684
rect 19180 47630 19182 47682
rect 19234 47630 19348 47682
rect 19180 47628 19348 47630
rect 19180 47618 19236 47628
rect 18956 47572 19012 47582
rect 19012 47516 19124 47572
rect 18956 47506 19012 47516
rect 18732 46946 18788 46956
rect 18844 47124 18900 47134
rect 18508 46834 18564 46844
rect 18732 46674 18788 46686
rect 18732 46622 18734 46674
rect 18786 46622 18788 46674
rect 18732 46452 18788 46622
rect 18844 46676 18900 47068
rect 18956 46676 19012 46686
rect 18844 46674 19012 46676
rect 18844 46622 18958 46674
rect 19010 46622 19012 46674
rect 18844 46620 19012 46622
rect 18956 46610 19012 46620
rect 18732 46386 18788 46396
rect 18732 46116 18788 46126
rect 18732 46002 18788 46060
rect 18732 45950 18734 46002
rect 18786 45950 18788 46002
rect 18732 45938 18788 45950
rect 18956 45892 19012 45902
rect 18956 45798 19012 45836
rect 19068 45892 19124 47516
rect 19292 47458 19348 47470
rect 19292 47406 19294 47458
rect 19346 47406 19348 47458
rect 19180 45892 19236 45902
rect 19068 45890 19236 45892
rect 19068 45838 19182 45890
rect 19234 45838 19236 45890
rect 19068 45836 19236 45838
rect 19068 45668 19124 45836
rect 19180 45826 19236 45836
rect 19292 45780 19348 47406
rect 19404 47348 19460 48412
rect 19404 47282 19460 47292
rect 19516 47684 19572 47694
rect 19404 46900 19460 46910
rect 19404 46450 19460 46844
rect 19404 46398 19406 46450
rect 19458 46398 19460 46450
rect 19404 46386 19460 46398
rect 19404 45780 19460 45790
rect 19292 45724 19404 45780
rect 19404 45714 19460 45724
rect 18732 45612 19124 45668
rect 19180 45668 19236 45678
rect 18732 45330 18788 45612
rect 18732 45278 18734 45330
rect 18786 45278 18788 45330
rect 18732 45266 18788 45278
rect 19068 44994 19124 45006
rect 19068 44942 19070 44994
rect 19122 44942 19124 44994
rect 19068 44884 19124 44942
rect 18956 44828 19068 44884
rect 18844 44436 18900 44446
rect 18844 44342 18900 44380
rect 18284 43820 18452 43876
rect 18508 44322 18564 44334
rect 18508 44270 18510 44322
rect 18562 44270 18564 44322
rect 18172 43540 18228 43550
rect 18060 43538 18228 43540
rect 18060 43486 18174 43538
rect 18226 43486 18228 43538
rect 18060 43484 18228 43486
rect 18060 42868 18116 43484
rect 18172 43474 18228 43484
rect 18284 43092 18340 43820
rect 18396 43650 18452 43662
rect 18396 43598 18398 43650
rect 18450 43598 18452 43650
rect 18396 43540 18452 43598
rect 18396 43474 18452 43484
rect 18060 42802 18116 42812
rect 18172 43036 18340 43092
rect 17836 41570 17892 41580
rect 17948 41858 18004 41870
rect 17948 41806 17950 41858
rect 18002 41806 18004 41858
rect 17948 41412 18004 41806
rect 17948 41346 18004 41356
rect 17948 41188 18004 41198
rect 18172 41188 18228 43036
rect 18508 42980 18564 44270
rect 18956 43876 19012 44828
rect 19068 44818 19124 44828
rect 18956 43810 19012 43820
rect 19068 44324 19124 44334
rect 19180 44324 19236 45612
rect 19516 45220 19572 47628
rect 19628 45332 19684 50316
rect 19964 50372 20020 50410
rect 20524 50372 20692 50428
rect 20748 50418 20804 50428
rect 19964 50306 20020 50316
rect 20524 50260 20580 50270
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 20188 49924 20244 49934
rect 20188 49830 20244 49868
rect 19852 49810 19908 49822
rect 19852 49758 19854 49810
rect 19906 49758 19908 49810
rect 19852 49476 19908 49758
rect 20412 49812 20468 49822
rect 19964 49700 20020 49710
rect 19964 49606 20020 49644
rect 19852 49410 19908 49420
rect 20188 49140 20244 49150
rect 20188 49046 20244 49084
rect 19964 49028 20020 49038
rect 19964 48934 20020 48972
rect 20300 48692 20356 48702
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 20188 48636 20300 48692
rect 20076 48244 20132 48254
rect 20076 48150 20132 48188
rect 20188 48132 20244 48636
rect 20300 48626 20356 48636
rect 19852 47684 19908 47694
rect 19852 47570 19908 47628
rect 19852 47518 19854 47570
rect 19906 47518 19908 47570
rect 19852 47506 19908 47518
rect 20188 47458 20244 48076
rect 20188 47406 20190 47458
rect 20242 47406 20244 47458
rect 20188 47394 20244 47406
rect 20300 47684 20356 47694
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 20300 46900 20356 47628
rect 20412 47236 20468 49756
rect 20412 47170 20468 47180
rect 20412 46900 20468 46910
rect 20300 46898 20468 46900
rect 20300 46846 20414 46898
rect 20466 46846 20468 46898
rect 20300 46844 20468 46846
rect 20412 46834 20468 46844
rect 19740 46674 19796 46686
rect 19740 46622 19742 46674
rect 19794 46622 19796 46674
rect 19740 46116 19796 46622
rect 20188 46674 20244 46686
rect 20188 46622 20190 46674
rect 20242 46622 20244 46674
rect 20188 46452 20244 46622
rect 20188 46386 20244 46396
rect 20300 46562 20356 46574
rect 20300 46510 20302 46562
rect 20354 46510 20356 46562
rect 20300 46228 20356 46510
rect 20300 46162 20356 46172
rect 19740 46050 19796 46060
rect 20412 46116 20468 46126
rect 20300 46004 20356 46014
rect 20412 46004 20468 46060
rect 20300 46002 20468 46004
rect 20300 45950 20302 46002
rect 20354 45950 20468 46002
rect 20300 45948 20468 45950
rect 20300 45938 20356 45948
rect 19740 45780 19796 45790
rect 19740 45686 19796 45724
rect 20188 45778 20244 45790
rect 20524 45780 20580 50204
rect 20636 49028 20692 50372
rect 20636 48962 20692 48972
rect 20636 48020 20692 48030
rect 20636 47926 20692 47964
rect 20748 47572 20804 47582
rect 20748 47478 20804 47516
rect 20748 47236 20804 47246
rect 20188 45726 20190 45778
rect 20242 45726 20244 45778
rect 20076 45668 20132 45678
rect 20188 45668 20244 45726
rect 20132 45612 20244 45668
rect 20412 45778 20580 45780
rect 20412 45726 20526 45778
rect 20578 45726 20580 45778
rect 20412 45724 20580 45726
rect 20076 45602 20132 45612
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 19628 45266 19684 45276
rect 19404 45164 19572 45220
rect 19740 45220 19796 45230
rect 19796 45164 19908 45220
rect 19292 44772 19348 44782
rect 19292 44546 19348 44716
rect 19292 44494 19294 44546
rect 19346 44494 19348 44546
rect 19292 44482 19348 44494
rect 19068 44322 19236 44324
rect 19068 44270 19070 44322
rect 19122 44270 19236 44322
rect 19068 44268 19236 44270
rect 18956 43538 19012 43550
rect 18956 43486 18958 43538
rect 19010 43486 19012 43538
rect 18284 42924 18564 42980
rect 18732 42980 18788 42990
rect 18284 42868 18340 42924
rect 18732 42886 18788 42924
rect 18284 42774 18340 42812
rect 18732 42756 18788 42766
rect 18732 42662 18788 42700
rect 18956 42084 19012 43486
rect 18956 42018 19012 42028
rect 18284 41970 18340 41982
rect 18284 41918 18286 41970
rect 18338 41918 18340 41970
rect 18284 41300 18340 41918
rect 18284 41234 18340 41244
rect 18396 41860 18452 41870
rect 18396 41746 18452 41804
rect 18396 41694 18398 41746
rect 18450 41694 18452 41746
rect 17948 41186 18228 41188
rect 17948 41134 17950 41186
rect 18002 41134 18174 41186
rect 18226 41134 18228 41186
rect 17948 41132 18228 41134
rect 17948 41122 18004 41132
rect 17164 38098 17220 38108
rect 17388 38612 17668 38668
rect 17724 41076 17780 41086
rect 17724 40516 17780 41020
rect 16268 37986 16324 37996
rect 16604 38050 16660 38062
rect 16604 37998 16606 38050
rect 16658 37998 16660 38050
rect 14028 37884 14756 37940
rect 15484 37828 15540 37838
rect 15596 37828 15652 37838
rect 15540 37826 15652 37828
rect 15540 37774 15598 37826
rect 15650 37774 15652 37826
rect 15540 37772 15652 37774
rect 14028 37380 14084 37390
rect 13692 37324 14028 37380
rect 14028 37286 14084 37324
rect 15148 37380 15204 37390
rect 15148 37286 15204 37324
rect 13132 37266 13188 37278
rect 13132 37214 13134 37266
rect 13186 37214 13188 37266
rect 13132 36708 13188 37214
rect 13580 37268 13636 37278
rect 13580 37266 13748 37268
rect 13580 37214 13582 37266
rect 13634 37214 13748 37266
rect 13580 37212 13748 37214
rect 13580 37202 13636 37212
rect 13132 36642 13188 36652
rect 13468 36596 13524 36606
rect 13468 36482 13524 36540
rect 13468 36430 13470 36482
rect 13522 36430 13524 36482
rect 13468 36418 13524 36430
rect 13580 36484 13636 36494
rect 12908 36318 12910 36370
rect 12962 36318 12964 36370
rect 12908 36260 12964 36318
rect 10668 35810 10836 35812
rect 10668 35758 10670 35810
rect 10722 35758 10836 35810
rect 10668 35756 10836 35758
rect 10668 35746 10724 35756
rect 11116 35700 11172 35710
rect 11116 35606 11172 35644
rect 11676 35700 11732 35710
rect 11900 35700 11956 36204
rect 12908 36194 12964 36204
rect 13580 35812 13636 36428
rect 13580 35718 13636 35756
rect 13692 36482 13748 37212
rect 15372 37266 15428 37278
rect 15372 37214 15374 37266
rect 15426 37214 15428 37266
rect 14588 36932 14644 36942
rect 15372 36932 15428 37214
rect 13692 36430 13694 36482
rect 13746 36430 13748 36482
rect 11676 35698 11900 35700
rect 11676 35646 11678 35698
rect 11730 35646 11900 35698
rect 11676 35644 11900 35646
rect 11676 35634 11732 35644
rect 11900 35606 11956 35644
rect 12012 35698 12068 35710
rect 12012 35646 12014 35698
rect 12066 35646 12068 35698
rect 12012 35364 12068 35646
rect 13244 35700 13300 35710
rect 13244 35606 13300 35644
rect 13692 35700 13748 36430
rect 13692 35634 13748 35644
rect 13916 36708 13972 36718
rect 12460 35588 12516 35598
rect 12460 35494 12516 35532
rect 12012 35298 12068 35308
rect 12908 35028 12964 35038
rect 12908 34934 12964 34972
rect 13468 35028 13524 35038
rect 13468 34914 13524 34972
rect 13468 34862 13470 34914
rect 13522 34862 13524 34914
rect 13468 34850 13524 34862
rect 10444 34750 10446 34802
rect 10498 34750 10500 34802
rect 9772 34692 9828 34702
rect 10108 34692 10164 34702
rect 9772 34690 10164 34692
rect 9772 34638 9774 34690
rect 9826 34638 10110 34690
rect 10162 34638 10164 34690
rect 9772 34636 10164 34638
rect 10444 34692 10500 34750
rect 11116 34804 11172 34814
rect 10892 34692 10948 34702
rect 10444 34690 10948 34692
rect 10444 34638 10894 34690
rect 10946 34638 10948 34690
rect 10444 34636 10948 34638
rect 9772 34626 9828 34636
rect 9100 34354 9716 34356
rect 9100 34302 9102 34354
rect 9154 34302 9716 34354
rect 9100 34300 9716 34302
rect 9996 34356 10052 34366
rect 9100 34290 9156 34300
rect 8988 34066 9044 34076
rect 9548 34130 9604 34142
rect 9548 34078 9550 34130
rect 9602 34078 9604 34130
rect 8540 33182 8542 33234
rect 8594 33182 8596 33234
rect 8540 33170 8596 33182
rect 9548 34020 9604 34078
rect 9100 33124 9156 33134
rect 9548 33124 9604 33964
rect 9996 34018 10052 34300
rect 9996 33966 9998 34018
rect 10050 33966 10052 34018
rect 9996 33954 10052 33966
rect 9100 33122 9604 33124
rect 9100 33070 9102 33122
rect 9154 33070 9604 33122
rect 9100 33068 9604 33070
rect 8428 32172 8820 32228
rect 7868 31166 7870 31218
rect 7922 31166 7924 31218
rect 5628 30046 5630 30098
rect 5682 30046 5684 30098
rect 5628 30034 5684 30046
rect 5964 30100 6020 30110
rect 5964 30006 6020 30044
rect 7868 30100 7924 31166
rect 8764 31218 8820 32172
rect 8764 31166 8766 31218
rect 8818 31166 8820 31218
rect 7868 30034 7924 30044
rect 8428 30770 8484 30782
rect 8428 30718 8430 30770
rect 8482 30718 8484 30770
rect 7756 29986 7812 29998
rect 7756 29934 7758 29986
rect 7810 29934 7812 29986
rect 7196 29876 7252 29886
rect 4620 27858 4900 27860
rect 4620 27806 4622 27858
rect 4674 27806 4900 27858
rect 4620 27804 4900 27806
rect 5068 29092 5124 29102
rect 5068 27858 5124 29036
rect 5068 27806 5070 27858
rect 5122 27806 5124 27858
rect 4620 27794 4676 27804
rect 5068 27794 5124 27806
rect 5964 28756 6020 28766
rect 1932 27636 1988 27646
rect 1932 27298 1988 27580
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 1932 27246 1934 27298
rect 1986 27246 1988 27298
rect 1932 27234 1988 27246
rect 4284 27074 4340 27086
rect 4284 27022 4286 27074
rect 4338 27022 4340 27074
rect 1708 26964 1764 26974
rect 1708 26514 1764 26908
rect 4284 26908 4340 27022
rect 4844 26964 4900 26974
rect 4284 26852 4900 26908
rect 1708 26462 1710 26514
rect 1762 26462 1764 26514
rect 1708 26450 1764 26462
rect 4844 26290 4900 26852
rect 4844 26238 4846 26290
rect 4898 26238 4900 26290
rect 4844 26226 4900 26238
rect 5068 26402 5124 26414
rect 5068 26350 5070 26402
rect 5122 26350 5124 26402
rect 2156 26066 2212 26078
rect 2156 26014 2158 26066
rect 2210 26014 2212 26066
rect 2156 25620 2212 26014
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 2156 25554 2212 25564
rect 1708 24500 1764 24510
rect 1708 24406 1764 24444
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 5068 23156 5124 26350
rect 5964 26178 6020 28700
rect 6972 28644 7028 28654
rect 6972 28550 7028 28588
rect 6636 28532 6692 28542
rect 6076 27076 6132 27086
rect 6076 26402 6132 27020
rect 6636 27074 6692 28476
rect 7196 28084 7252 29820
rect 7756 28756 7812 29934
rect 7756 28690 7812 28700
rect 7644 28644 7700 28654
rect 7308 28420 7364 28430
rect 7308 28418 7588 28420
rect 7308 28366 7310 28418
rect 7362 28366 7588 28418
rect 7308 28364 7588 28366
rect 7308 28354 7364 28364
rect 7308 28084 7364 28094
rect 7196 28082 7364 28084
rect 7196 28030 7310 28082
rect 7362 28030 7364 28082
rect 7196 28028 7364 28030
rect 7308 28018 7364 28028
rect 6636 27022 6638 27074
rect 6690 27022 6692 27074
rect 6636 27010 6692 27022
rect 7308 27636 7364 27646
rect 7308 27076 7364 27580
rect 7308 26982 7364 27020
rect 7532 27076 7588 28364
rect 7644 27188 7700 28588
rect 8428 28532 8484 30718
rect 8764 30212 8820 31166
rect 8540 30100 8596 30110
rect 8540 30006 8596 30044
rect 8428 27972 8484 28476
rect 8764 28084 8820 30156
rect 9100 29876 9156 33068
rect 10108 31780 10164 34636
rect 10556 34468 10612 34478
rect 10556 34354 10612 34412
rect 10556 34302 10558 34354
rect 10610 34302 10612 34354
rect 10556 34290 10612 34302
rect 10892 32788 10948 34636
rect 11116 34354 11172 34748
rect 13804 34804 13860 34814
rect 13916 34804 13972 36652
rect 14588 36706 14644 36876
rect 15260 36876 15372 36932
rect 14588 36654 14590 36706
rect 14642 36654 14644 36706
rect 14588 36642 14644 36654
rect 14924 36708 14980 36718
rect 14140 36482 14196 36494
rect 14140 36430 14142 36482
rect 14194 36430 14196 36482
rect 14140 36148 14196 36430
rect 14140 35700 14196 36092
rect 14252 35924 14308 35934
rect 14252 35830 14308 35868
rect 14924 35810 14980 36652
rect 15260 36596 15316 36876
rect 15372 36866 15428 36876
rect 14924 35758 14926 35810
rect 14978 35758 14980 35810
rect 14140 35606 14196 35644
rect 14812 35700 14868 35710
rect 14812 35606 14868 35644
rect 13804 34802 13972 34804
rect 13804 34750 13806 34802
rect 13858 34750 13972 34802
rect 13804 34748 13972 34750
rect 14028 35252 14084 35262
rect 13804 34738 13860 34748
rect 11340 34692 11396 34702
rect 11340 34598 11396 34636
rect 11116 34302 11118 34354
rect 11170 34302 11172 34354
rect 11116 33684 11172 34302
rect 13692 34130 13748 34142
rect 13692 34078 13694 34130
rect 13746 34078 13748 34130
rect 11116 33618 11172 33628
rect 13020 33684 13076 33694
rect 11676 33348 11732 33358
rect 11676 33254 11732 33292
rect 12012 33346 12068 33358
rect 12012 33294 12014 33346
rect 12066 33294 12068 33346
rect 10892 32722 10948 32732
rect 12012 33124 12068 33294
rect 10108 31714 10164 31724
rect 11788 32452 11844 32462
rect 12012 32452 12068 33068
rect 12572 33124 12628 33134
rect 12572 33030 12628 33068
rect 11788 32450 12068 32452
rect 11788 32398 11790 32450
rect 11842 32398 12068 32450
rect 11788 32396 12068 32398
rect 9884 31106 9940 31118
rect 9884 31054 9886 31106
rect 9938 31054 9940 31106
rect 9660 30996 9716 31006
rect 9660 30994 9828 30996
rect 9660 30942 9662 30994
rect 9714 30942 9828 30994
rect 9660 30940 9828 30942
rect 9660 30930 9716 30940
rect 9772 29876 9828 30940
rect 9884 30100 9940 31054
rect 9884 30034 9940 30044
rect 10780 30210 10836 30222
rect 10780 30158 10782 30210
rect 10834 30158 10836 30210
rect 10780 30100 10836 30158
rect 11228 30212 11284 30222
rect 11228 30118 11284 30156
rect 11788 30212 11844 32396
rect 13020 31218 13076 33628
rect 13692 33236 13748 34078
rect 14028 33570 14084 35196
rect 14476 35028 14532 35038
rect 14252 34690 14308 34702
rect 14252 34638 14254 34690
rect 14306 34638 14308 34690
rect 14252 34468 14308 34638
rect 14252 34402 14308 34412
rect 14476 34354 14532 34972
rect 14812 34916 14868 34926
rect 14924 34916 14980 35758
rect 14812 34914 14980 34916
rect 14812 34862 14814 34914
rect 14866 34862 14980 34914
rect 14812 34860 14980 34862
rect 15036 36540 15316 36596
rect 14812 34850 14868 34860
rect 15036 34802 15092 36540
rect 15484 36482 15540 37772
rect 15596 37762 15652 37772
rect 15932 37492 15988 37502
rect 15932 37398 15988 37436
rect 15596 37268 15652 37278
rect 15596 36932 15652 37212
rect 16604 36932 16660 37998
rect 15596 36876 16212 36932
rect 15484 36430 15486 36482
rect 15538 36430 15540 36482
rect 15372 36370 15428 36382
rect 15372 36318 15374 36370
rect 15426 36318 15428 36370
rect 15372 35812 15428 36318
rect 15484 36036 15540 36430
rect 15708 36370 15764 36382
rect 15708 36318 15710 36370
rect 15762 36318 15764 36370
rect 15708 36148 15764 36318
rect 16156 36370 16212 36876
rect 16156 36318 16158 36370
rect 16210 36318 16212 36370
rect 16156 36306 16212 36318
rect 16380 36482 16436 36494
rect 16380 36430 16382 36482
rect 16434 36430 16436 36482
rect 16380 36148 16436 36430
rect 16604 36484 16660 36876
rect 17164 36484 17220 36494
rect 16604 36482 17220 36484
rect 16604 36430 17166 36482
rect 17218 36430 17220 36482
rect 16604 36428 17220 36430
rect 15708 36092 16436 36148
rect 15484 35980 15988 36036
rect 15708 35812 15764 35822
rect 15428 35810 15764 35812
rect 15428 35758 15710 35810
rect 15762 35758 15764 35810
rect 15428 35756 15764 35758
rect 15372 35718 15428 35756
rect 15708 35746 15764 35756
rect 15932 35698 15988 35980
rect 16268 35924 16324 35934
rect 16268 35830 16324 35868
rect 15932 35646 15934 35698
rect 15986 35646 15988 35698
rect 15932 35634 15988 35646
rect 15372 35586 15428 35598
rect 15372 35534 15374 35586
rect 15426 35534 15428 35586
rect 15372 34916 15428 35534
rect 15372 34850 15428 34860
rect 15036 34750 15038 34802
rect 15090 34750 15092 34802
rect 15036 34738 15092 34750
rect 16380 34804 16436 36092
rect 17052 36258 17108 36270
rect 17052 36206 17054 36258
rect 17106 36206 17108 36258
rect 17052 36148 17108 36206
rect 17052 36082 17108 36092
rect 17164 35924 17220 36428
rect 17388 36148 17444 38612
rect 17388 36082 17444 36092
rect 17500 38500 17556 38510
rect 17388 35924 17444 35934
rect 17164 35922 17444 35924
rect 17164 35870 17390 35922
rect 17442 35870 17444 35922
rect 17164 35868 17444 35870
rect 17388 35858 17444 35868
rect 17500 35812 17556 38444
rect 17612 37492 17668 37502
rect 17612 37398 17668 37436
rect 17724 36484 17780 40460
rect 17836 40402 17892 40414
rect 17836 40350 17838 40402
rect 17890 40350 17892 40402
rect 17836 40292 17892 40350
rect 17836 39508 17892 40236
rect 17836 38946 17892 39452
rect 17836 38894 17838 38946
rect 17890 38894 17892 38946
rect 17836 38882 17892 38894
rect 17948 39620 18004 39630
rect 17948 38836 18004 39564
rect 17948 38742 18004 38780
rect 17836 38052 17892 38062
rect 17836 37958 17892 37996
rect 17948 37828 18004 37838
rect 17948 37154 18004 37772
rect 18172 37268 18228 41132
rect 18396 41188 18452 41694
rect 18396 41122 18452 41132
rect 18844 41298 18900 41310
rect 18844 41246 18846 41298
rect 18898 41246 18900 41298
rect 18844 40852 18900 41246
rect 18956 41300 19012 41310
rect 18956 41186 19012 41244
rect 18956 41134 18958 41186
rect 19010 41134 19012 41186
rect 18956 41122 19012 41134
rect 19068 40852 19124 44268
rect 19404 43652 19460 45164
rect 19740 45154 19796 45164
rect 19852 45106 19908 45164
rect 19852 45054 19854 45106
rect 19906 45054 19908 45106
rect 19516 44996 19572 45006
rect 19852 44996 19908 45054
rect 19516 44994 19908 44996
rect 19516 44942 19518 44994
rect 19570 44942 19908 44994
rect 19516 44940 19908 44942
rect 19964 45218 20020 45230
rect 19964 45166 19966 45218
rect 20018 45166 20020 45218
rect 19964 45108 20020 45166
rect 20188 45220 20244 45230
rect 20188 45126 20244 45164
rect 19516 44930 19572 44940
rect 19964 44660 20020 45052
rect 19852 44604 20020 44660
rect 19404 43586 19460 43596
rect 19516 44548 19572 44558
rect 19516 44324 19572 44492
rect 19516 43538 19572 44268
rect 19852 44324 19908 44604
rect 19852 44230 19908 44268
rect 19964 44212 20020 44222
rect 19964 44118 20020 44156
rect 20188 44098 20244 44110
rect 20188 44046 20190 44098
rect 20242 44046 20244 44098
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 19740 43652 19796 43662
rect 19796 43596 19908 43652
rect 19740 43586 19796 43596
rect 19516 43486 19518 43538
rect 19570 43486 19572 43538
rect 19516 43474 19572 43486
rect 19740 43428 19796 43438
rect 19516 42868 19572 42878
rect 18844 40786 18900 40796
rect 18956 40796 19124 40852
rect 19180 42866 19572 42868
rect 19180 42814 19518 42866
rect 19570 42814 19572 42866
rect 19180 42812 19572 42814
rect 18956 40292 19012 40796
rect 19180 40628 19236 42812
rect 19516 42802 19572 42812
rect 19740 42754 19796 43372
rect 19740 42702 19742 42754
rect 19794 42702 19796 42754
rect 19740 42690 19796 42702
rect 19404 42644 19460 42654
rect 19404 42550 19460 42588
rect 19852 42532 19908 43596
rect 20188 43540 20244 44046
rect 20412 43876 20468 45724
rect 20524 45714 20580 45724
rect 20636 46450 20692 46462
rect 20636 46398 20638 46450
rect 20690 46398 20692 46450
rect 20524 45108 20580 45118
rect 20636 45108 20692 46398
rect 20524 45106 20692 45108
rect 20524 45054 20526 45106
rect 20578 45054 20692 45106
rect 20524 45052 20692 45054
rect 20748 45778 20804 47180
rect 20860 46004 20916 51326
rect 20972 49028 21028 56140
rect 21868 56196 21924 56206
rect 21868 56102 21924 56140
rect 22652 56196 22708 56206
rect 21308 56084 21364 56094
rect 21308 55990 21364 56028
rect 21756 55860 21812 55870
rect 21756 55298 21812 55804
rect 22540 55636 22596 55646
rect 22652 55636 22708 56140
rect 22596 55580 22708 55636
rect 22540 55570 22596 55580
rect 21756 55246 21758 55298
rect 21810 55246 21812 55298
rect 21196 54626 21252 54638
rect 21196 54574 21198 54626
rect 21250 54574 21252 54626
rect 21196 53956 21252 54574
rect 21756 54628 21812 55246
rect 22428 55412 22484 55422
rect 22204 55188 22260 55198
rect 22204 55094 22260 55132
rect 21756 54562 21812 54572
rect 22428 54516 22484 55356
rect 22652 55410 22708 55580
rect 22652 55358 22654 55410
rect 22706 55358 22708 55410
rect 22652 55346 22708 55358
rect 22764 55636 22820 55646
rect 22652 54740 22708 54750
rect 22652 54646 22708 54684
rect 22428 54514 22596 54516
rect 22428 54462 22430 54514
rect 22482 54462 22596 54514
rect 22428 54460 22596 54462
rect 22428 54450 22484 54460
rect 22092 54292 22148 54302
rect 21196 53890 21252 53900
rect 21980 54236 22092 54292
rect 21532 53732 21588 53742
rect 21532 53730 21700 53732
rect 21532 53678 21534 53730
rect 21586 53678 21700 53730
rect 21532 53676 21700 53678
rect 21532 53666 21588 53676
rect 21308 52948 21364 52958
rect 21308 52854 21364 52892
rect 21644 52836 21700 53676
rect 21420 52500 21476 52510
rect 21420 52276 21476 52444
rect 21084 52164 21140 52174
rect 21084 50484 21140 52108
rect 21420 52162 21476 52220
rect 21420 52110 21422 52162
rect 21474 52110 21476 52162
rect 21420 52098 21476 52110
rect 21644 52164 21700 52780
rect 21644 52098 21700 52108
rect 21532 52050 21588 52062
rect 21532 51998 21534 52050
rect 21586 51998 21588 52050
rect 21532 51940 21588 51998
rect 21420 51884 21588 51940
rect 21196 51828 21252 51838
rect 21196 51380 21252 51772
rect 21196 51286 21252 51324
rect 21420 51156 21476 51884
rect 21868 51604 21924 51614
rect 21756 51492 21812 51502
rect 21084 50418 21140 50428
rect 21196 51100 21476 51156
rect 21532 51378 21588 51390
rect 21532 51326 21534 51378
rect 21586 51326 21588 51378
rect 21196 50708 21252 51100
rect 20972 48962 21028 48972
rect 21084 49924 21140 49934
rect 21084 48242 21140 49868
rect 21084 48190 21086 48242
rect 21138 48190 21140 48242
rect 20972 47124 21028 47134
rect 20972 46898 21028 47068
rect 20972 46846 20974 46898
rect 21026 46846 21028 46898
rect 20972 46834 21028 46846
rect 21084 46788 21140 48190
rect 21196 47236 21252 50652
rect 21308 50594 21364 50606
rect 21308 50542 21310 50594
rect 21362 50542 21364 50594
rect 21308 49588 21364 50542
rect 21420 50372 21476 50382
rect 21420 49922 21476 50316
rect 21420 49870 21422 49922
rect 21474 49870 21476 49922
rect 21420 49858 21476 49870
rect 21308 49522 21364 49532
rect 21308 49028 21364 49038
rect 21308 47458 21364 48972
rect 21308 47406 21310 47458
rect 21362 47406 21364 47458
rect 21308 47394 21364 47406
rect 21420 47348 21476 47358
rect 21532 47348 21588 51326
rect 21644 51268 21700 51278
rect 21644 50594 21700 51212
rect 21644 50542 21646 50594
rect 21698 50542 21700 50594
rect 21644 50530 21700 50542
rect 21644 50372 21700 50382
rect 21644 49810 21700 50316
rect 21644 49758 21646 49810
rect 21698 49758 21700 49810
rect 21644 49746 21700 49758
rect 21644 49588 21700 49598
rect 21644 47684 21700 49532
rect 21756 49026 21812 51436
rect 21756 48974 21758 49026
rect 21810 48974 21812 49026
rect 21756 48962 21812 48974
rect 21644 47618 21700 47628
rect 21756 48244 21812 48254
rect 21420 47346 21588 47348
rect 21420 47294 21422 47346
rect 21474 47294 21588 47346
rect 21420 47292 21588 47294
rect 21196 47180 21364 47236
rect 21084 46722 21140 46732
rect 21308 46786 21364 47180
rect 21308 46734 21310 46786
rect 21362 46734 21364 46786
rect 21308 46676 21364 46734
rect 21196 46620 21364 46676
rect 21196 46564 21252 46620
rect 21420 46564 21476 47292
rect 21084 46508 21252 46564
rect 21308 46508 21476 46564
rect 21084 46450 21140 46508
rect 21308 46452 21364 46508
rect 21532 46452 21588 46462
rect 21084 46398 21086 46450
rect 21138 46398 21140 46450
rect 21084 46386 21140 46398
rect 21196 46396 21364 46452
rect 21420 46450 21588 46452
rect 21420 46398 21534 46450
rect 21586 46398 21588 46450
rect 21420 46396 21588 46398
rect 20860 45938 20916 45948
rect 20748 45726 20750 45778
rect 20802 45726 20804 45778
rect 20748 45218 20804 45726
rect 20748 45166 20750 45218
rect 20802 45166 20804 45218
rect 20524 45042 20580 45052
rect 20524 44884 20580 44894
rect 20580 44828 20692 44884
rect 20524 44818 20580 44828
rect 20524 44212 20580 44222
rect 20524 44118 20580 44156
rect 20412 43820 20580 43876
rect 20412 43652 20468 43662
rect 20412 43540 20468 43596
rect 20188 43538 20468 43540
rect 20188 43486 20414 43538
rect 20466 43486 20468 43538
rect 20188 43484 20468 43486
rect 20412 43474 20468 43484
rect 20412 42980 20468 42990
rect 20524 42980 20580 43820
rect 20468 42924 20580 42980
rect 20412 42914 20468 42924
rect 20524 42756 20580 42766
rect 20636 42756 20692 44828
rect 20748 44100 20804 45166
rect 20748 44034 20804 44044
rect 20972 45556 21028 45566
rect 20972 43538 21028 45500
rect 21196 44996 21252 46396
rect 21308 46116 21364 46126
rect 21308 45890 21364 46060
rect 21308 45838 21310 45890
rect 21362 45838 21364 45890
rect 21308 45826 21364 45838
rect 21196 44902 21252 44940
rect 21308 44324 21364 44334
rect 21308 44230 21364 44268
rect 21084 43652 21140 43662
rect 21084 43558 21140 43596
rect 20972 43486 20974 43538
rect 21026 43486 21028 43538
rect 20860 43316 20916 43326
rect 20524 42754 20692 42756
rect 20524 42702 20526 42754
rect 20578 42702 20692 42754
rect 20524 42700 20692 42702
rect 20748 43260 20860 43316
rect 20524 42690 20580 42700
rect 19628 42476 19908 42532
rect 19292 42084 19348 42094
rect 19292 41636 19348 42028
rect 19628 42082 19684 42476
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20748 42308 20804 43260
rect 20860 43250 20916 43260
rect 19836 42298 20100 42308
rect 20636 42252 20804 42308
rect 20860 42868 20916 42878
rect 19628 42030 19630 42082
rect 19682 42030 19684 42082
rect 19628 42018 19684 42030
rect 19964 42084 20020 42094
rect 19964 41990 20020 42028
rect 19404 41972 19460 41982
rect 19404 41878 19460 41916
rect 19740 41972 19796 41982
rect 19292 41580 19460 41636
rect 19292 41412 19348 41422
rect 19292 41076 19348 41356
rect 19292 41010 19348 41020
rect 18956 39956 19012 40236
rect 18956 39890 19012 39900
rect 19068 40572 19236 40628
rect 18396 39732 18452 39742
rect 18284 39396 18340 39406
rect 18284 38834 18340 39340
rect 18396 39058 18452 39676
rect 18396 39006 18398 39058
rect 18450 39006 18452 39058
rect 18396 38994 18452 39006
rect 18956 39396 19012 39406
rect 18284 38782 18286 38834
rect 18338 38782 18340 38834
rect 18284 38668 18340 38782
rect 18284 38612 18788 38668
rect 18732 38050 18788 38612
rect 18732 37998 18734 38050
rect 18786 37998 18788 38050
rect 18732 37986 18788 37998
rect 18396 37940 18452 37950
rect 18508 37940 18564 37950
rect 18396 37938 18508 37940
rect 18396 37886 18398 37938
rect 18450 37886 18508 37938
rect 18396 37884 18508 37886
rect 18396 37874 18452 37884
rect 18284 37268 18340 37278
rect 18172 37266 18340 37268
rect 18172 37214 18286 37266
rect 18338 37214 18340 37266
rect 18172 37212 18340 37214
rect 17948 37102 17950 37154
rect 18002 37102 18004 37154
rect 17948 37090 18004 37102
rect 17500 35746 17556 35756
rect 17612 36428 17780 36484
rect 18284 36820 18340 37212
rect 17612 35588 17668 36428
rect 17724 36260 17780 36270
rect 18060 36260 18116 36270
rect 17780 36258 18116 36260
rect 17780 36206 18062 36258
rect 18114 36206 18116 36258
rect 17780 36204 18116 36206
rect 17724 36166 17780 36204
rect 18060 36194 18116 36204
rect 17836 35588 17892 35598
rect 17612 35586 17892 35588
rect 17612 35534 17838 35586
rect 17890 35534 17892 35586
rect 17612 35532 17892 35534
rect 16380 34738 16436 34748
rect 16828 35252 16884 35262
rect 14476 34302 14478 34354
rect 14530 34302 14532 34354
rect 14476 34290 14532 34302
rect 14700 34468 14756 34478
rect 14028 33518 14030 33570
rect 14082 33518 14084 33570
rect 14028 33506 14084 33518
rect 14140 34130 14196 34142
rect 14140 34078 14142 34130
rect 14194 34078 14196 34130
rect 14140 34020 14196 34078
rect 14700 34130 14756 34412
rect 16828 34356 16884 35196
rect 17836 35028 17892 35532
rect 18284 35308 18340 36764
rect 18396 36372 18452 36382
rect 18396 36278 18452 36316
rect 18172 35252 18340 35308
rect 17836 34962 17892 34972
rect 18060 35028 18116 35038
rect 18172 35028 18228 35252
rect 18060 35026 18340 35028
rect 18060 34974 18062 35026
rect 18114 34974 18340 35026
rect 18060 34972 18340 34974
rect 18060 34962 18116 34972
rect 17388 34356 17444 34366
rect 16828 34354 17444 34356
rect 16828 34302 16830 34354
rect 16882 34302 17390 34354
rect 17442 34302 17444 34354
rect 16828 34300 17444 34302
rect 16828 34290 16884 34300
rect 17388 34290 17444 34300
rect 18284 34244 18340 34972
rect 18396 34804 18452 34814
rect 18396 34468 18452 34748
rect 18508 34580 18564 37884
rect 18732 37492 18788 37502
rect 18732 37398 18788 37436
rect 18956 37268 19012 39340
rect 19068 38612 19124 40572
rect 19180 40404 19236 40414
rect 19180 39730 19236 40348
rect 19180 39678 19182 39730
rect 19234 39678 19236 39730
rect 19180 39666 19236 39678
rect 19292 40402 19348 40414
rect 19292 40350 19294 40402
rect 19346 40350 19348 40402
rect 19292 39620 19348 40350
rect 19292 39526 19348 39564
rect 19180 39284 19236 39294
rect 19180 39058 19236 39228
rect 19180 39006 19182 39058
rect 19234 39006 19236 39058
rect 19180 38994 19236 39006
rect 19404 38948 19460 41580
rect 19628 41412 19684 41422
rect 19740 41412 19796 41916
rect 19684 41356 19796 41412
rect 20188 41636 20244 41646
rect 19628 41346 19684 41356
rect 19628 41076 19684 41086
rect 19628 40982 19684 41020
rect 20076 40964 20132 41002
rect 20076 40898 20132 40908
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19740 40628 19796 40638
rect 19740 40290 19796 40572
rect 19740 40238 19742 40290
rect 19794 40238 19796 40290
rect 19740 40226 19796 40238
rect 19740 39508 19796 39518
rect 19740 39414 19796 39452
rect 19516 39284 19572 39294
rect 19516 39058 19572 39228
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19516 39006 19518 39058
rect 19570 39006 19572 39058
rect 19516 38994 19572 39006
rect 19068 38546 19124 38556
rect 19292 38892 19460 38948
rect 19292 38388 19348 38892
rect 19964 38724 20020 38734
rect 19964 38630 20020 38668
rect 19068 38332 19348 38388
rect 19068 37492 19124 38332
rect 19292 38164 19348 38174
rect 19292 38070 19348 38108
rect 19628 38052 19684 38062
rect 19628 37828 19684 37996
rect 19740 37828 19796 37838
rect 19628 37826 19796 37828
rect 19628 37774 19742 37826
rect 19794 37774 19796 37826
rect 19628 37772 19796 37774
rect 19068 37490 19572 37492
rect 19068 37438 19070 37490
rect 19122 37438 19572 37490
rect 19068 37436 19572 37438
rect 19068 37426 19124 37436
rect 18956 37212 19124 37268
rect 18844 36820 18900 36830
rect 18844 36594 18900 36764
rect 18844 36542 18846 36594
rect 18898 36542 18900 36594
rect 18844 36530 18900 36542
rect 18956 36484 19012 36494
rect 18956 35308 19012 36428
rect 19068 35924 19124 37212
rect 19516 37156 19572 37436
rect 19628 37378 19684 37772
rect 19740 37762 19796 37772
rect 20188 37828 20244 41580
rect 20524 41076 20580 41086
rect 20188 37734 20244 37772
rect 20300 38612 20356 38622
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19628 37326 19630 37378
rect 19682 37326 19684 37378
rect 19628 37314 19684 37326
rect 19852 37266 19908 37278
rect 19852 37214 19854 37266
rect 19906 37214 19908 37266
rect 19852 37156 19908 37214
rect 19516 37100 19796 37156
rect 19404 36594 19460 36606
rect 19404 36542 19406 36594
rect 19458 36542 19460 36594
rect 19404 36484 19460 36542
rect 19404 36418 19460 36428
rect 19740 36482 19796 37100
rect 19740 36430 19742 36482
rect 19794 36430 19796 36482
rect 19740 36418 19796 36430
rect 19852 36260 19908 37100
rect 20188 37268 20244 37278
rect 20188 37154 20244 37212
rect 20188 37102 20190 37154
rect 20242 37102 20244 37154
rect 20188 37090 20244 37102
rect 20188 36596 20244 36606
rect 20300 36596 20356 38556
rect 20524 38276 20580 41020
rect 20636 39844 20692 42252
rect 20748 42082 20804 42094
rect 20748 42030 20750 42082
rect 20802 42030 20804 42082
rect 20748 41076 20804 42030
rect 20860 41298 20916 42812
rect 20860 41246 20862 41298
rect 20914 41246 20916 41298
rect 20860 41234 20916 41246
rect 20748 41010 20804 41020
rect 20748 40852 20804 40862
rect 20748 40628 20804 40796
rect 20748 40534 20804 40572
rect 20636 39778 20692 39788
rect 20748 40068 20804 40078
rect 20748 39730 20804 40012
rect 20748 39678 20750 39730
rect 20802 39678 20804 39730
rect 20748 39666 20804 39678
rect 20748 39284 20804 39294
rect 20748 39058 20804 39228
rect 20748 39006 20750 39058
rect 20802 39006 20804 39058
rect 20748 38994 20804 39006
rect 20860 38948 20916 38958
rect 20860 38854 20916 38892
rect 20636 38612 20692 38622
rect 20636 38518 20692 38556
rect 20412 38220 20580 38276
rect 20412 36932 20468 38220
rect 20748 38052 20804 38062
rect 20748 37958 20804 37996
rect 20524 37266 20580 37278
rect 20748 37268 20804 37278
rect 20524 37214 20526 37266
rect 20578 37214 20580 37266
rect 20524 37156 20580 37214
rect 20524 37090 20580 37100
rect 20636 37266 20804 37268
rect 20636 37214 20750 37266
rect 20802 37214 20804 37266
rect 20636 37212 20804 37214
rect 20412 36876 20580 36932
rect 20244 36540 20356 36596
rect 20188 36482 20244 36540
rect 20188 36430 20190 36482
rect 20242 36430 20244 36482
rect 20188 36418 20244 36430
rect 19628 36204 19908 36260
rect 19516 36148 19572 36158
rect 19068 35922 19460 35924
rect 19068 35870 19070 35922
rect 19122 35870 19460 35922
rect 19068 35868 19460 35870
rect 19068 35858 19124 35868
rect 18956 35252 19236 35308
rect 18732 35026 18788 35038
rect 18732 34974 18734 35026
rect 18786 34974 18788 35026
rect 18620 34916 18676 34926
rect 18620 34802 18676 34860
rect 18620 34750 18622 34802
rect 18674 34750 18676 34802
rect 18620 34738 18676 34750
rect 18508 34524 18676 34580
rect 18396 34412 18564 34468
rect 18396 34244 18452 34254
rect 14700 34078 14702 34130
rect 14754 34078 14756 34130
rect 14700 34066 14756 34078
rect 17948 34242 18452 34244
rect 17948 34190 18398 34242
rect 18450 34190 18452 34242
rect 17948 34188 18452 34190
rect 17948 34130 18004 34188
rect 18396 34178 18452 34188
rect 17948 34078 17950 34130
rect 18002 34078 18004 34130
rect 17948 34066 18004 34078
rect 13692 33170 13748 33180
rect 13580 33124 13636 33134
rect 13580 33030 13636 33068
rect 14028 33124 14084 33134
rect 14140 33124 14196 33964
rect 15260 34020 15316 34030
rect 14084 33068 14196 33124
rect 14588 33572 14644 33582
rect 14588 33122 14644 33516
rect 15260 33348 15316 33964
rect 18396 34020 18452 34030
rect 18508 34020 18564 34412
rect 18452 33964 18564 34020
rect 18396 33954 18452 33964
rect 18508 33796 18564 33806
rect 18620 33796 18676 34524
rect 18564 33740 18676 33796
rect 18732 34130 18788 34974
rect 19068 34468 19124 34478
rect 19068 34242 19124 34412
rect 19068 34190 19070 34242
rect 19122 34190 19124 34242
rect 19068 34178 19124 34190
rect 18732 34078 18734 34130
rect 18786 34078 18788 34130
rect 17164 33460 17220 33470
rect 15260 33282 15316 33292
rect 16604 33348 16660 33358
rect 14588 33070 14590 33122
rect 14642 33070 14644 33122
rect 14028 33058 14084 33068
rect 14588 33058 14644 33070
rect 16604 31220 16660 33292
rect 17164 33346 17220 33404
rect 18508 33458 18564 33740
rect 18732 33572 18788 34078
rect 19180 33908 19236 35252
rect 18732 33506 18788 33516
rect 18844 33852 19236 33908
rect 19292 35252 19348 35262
rect 18508 33406 18510 33458
rect 18562 33406 18564 33458
rect 18508 33394 18564 33406
rect 17164 33294 17166 33346
rect 17218 33294 17220 33346
rect 17164 33282 17220 33294
rect 17500 33348 17556 33358
rect 17500 33254 17556 33292
rect 18844 33346 18900 33852
rect 19292 33458 19348 35196
rect 19404 34916 19460 35868
rect 19404 34822 19460 34860
rect 19516 34356 19572 36092
rect 19628 35924 19684 36204
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19852 35924 19908 35934
rect 19628 35868 19852 35924
rect 19852 35830 19908 35868
rect 20412 35700 20468 35710
rect 20412 35606 20468 35644
rect 20076 35252 20132 35262
rect 20076 35138 20132 35196
rect 20076 35086 20078 35138
rect 20130 35086 20132 35138
rect 20076 35074 20132 35086
rect 19628 35028 19684 35038
rect 19628 34914 19684 34972
rect 19628 34862 19630 34914
rect 19682 34862 19684 34914
rect 19628 34850 19684 34862
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19516 34290 19572 34300
rect 19852 34356 19908 34366
rect 19628 34244 19684 34254
rect 19628 34150 19684 34188
rect 19516 34132 19572 34142
rect 19292 33406 19294 33458
rect 19346 33406 19348 33458
rect 19292 33394 19348 33406
rect 19404 34076 19516 34132
rect 18844 33294 18846 33346
rect 18898 33294 18900 33346
rect 18844 33282 18900 33294
rect 18956 33124 19012 33134
rect 18956 33030 19012 33068
rect 19068 33122 19124 33134
rect 19068 33070 19070 33122
rect 19122 33070 19124 33122
rect 18508 32676 18564 32686
rect 13020 31166 13022 31218
rect 13074 31166 13076 31218
rect 13020 31154 13076 31166
rect 16156 31218 16660 31220
rect 16156 31166 16606 31218
rect 16658 31166 16660 31218
rect 16156 31164 16660 31166
rect 15484 30994 15540 31006
rect 15484 30942 15486 30994
rect 15538 30942 15540 30994
rect 11788 30118 11844 30156
rect 12460 30770 12516 30782
rect 12460 30718 12462 30770
rect 12514 30718 12516 30770
rect 10780 30034 10836 30044
rect 9772 29820 10164 29876
rect 9100 29810 9156 29820
rect 10108 29538 10164 29820
rect 10108 29486 10110 29538
rect 10162 29486 10164 29538
rect 10108 29474 10164 29486
rect 10556 29428 10612 29438
rect 10444 29426 10612 29428
rect 10444 29374 10558 29426
rect 10610 29374 10612 29426
rect 10444 29372 10612 29374
rect 9772 29316 9828 29326
rect 9772 29222 9828 29260
rect 10444 29316 10500 29372
rect 10556 29362 10612 29372
rect 11004 29428 11060 29438
rect 11004 29334 11060 29372
rect 9212 28644 9268 28654
rect 9100 28420 9156 28430
rect 8988 28364 9100 28420
rect 8876 28084 8932 28094
rect 8764 28082 8932 28084
rect 8764 28030 8878 28082
rect 8930 28030 8932 28082
rect 8764 28028 8932 28030
rect 8876 28018 8932 28028
rect 8428 27878 8484 27916
rect 8092 27636 8148 27646
rect 8316 27636 8372 27646
rect 8988 27636 9044 28364
rect 9100 28354 9156 28364
rect 9212 28418 9268 28588
rect 9212 28366 9214 28418
rect 9266 28366 9268 28418
rect 8092 27542 8148 27580
rect 8204 27634 8372 27636
rect 8204 27582 8318 27634
rect 8370 27582 8372 27634
rect 8204 27580 8372 27582
rect 7644 27186 8148 27188
rect 7644 27134 7646 27186
rect 7698 27134 8148 27186
rect 7644 27132 8148 27134
rect 7644 27122 7700 27132
rect 6860 26852 6916 26862
rect 6860 26850 7140 26852
rect 6860 26798 6862 26850
rect 6914 26798 7140 26850
rect 6860 26796 7140 26798
rect 6860 26786 6916 26796
rect 6076 26350 6078 26402
rect 6130 26350 6132 26402
rect 6076 26338 6132 26350
rect 5964 26126 5966 26178
rect 6018 26126 6020 26178
rect 5964 26114 6020 26126
rect 6860 26180 6916 26190
rect 6860 26086 6916 26124
rect 6412 25844 6468 25854
rect 5964 25508 6020 25518
rect 5964 25414 6020 25452
rect 5628 25396 5684 25406
rect 5628 24050 5684 25340
rect 6076 24724 6132 24734
rect 5740 24722 6132 24724
rect 5740 24670 6078 24722
rect 6130 24670 6132 24722
rect 5740 24668 6132 24670
rect 5740 24162 5796 24668
rect 5740 24110 5742 24162
rect 5794 24110 5796 24162
rect 5740 24098 5796 24110
rect 5628 23998 5630 24050
rect 5682 23998 5684 24050
rect 5628 23156 5684 23998
rect 5068 23154 5348 23156
rect 5068 23102 5070 23154
rect 5122 23102 5348 23154
rect 5068 23100 5348 23102
rect 5068 23090 5124 23100
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 1708 21698 1764 21710
rect 1708 21646 1710 21698
rect 1762 21646 1764 21698
rect 1708 20916 1764 21646
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 1708 20850 1764 20860
rect 5292 20132 5348 23100
rect 5628 23154 5908 23156
rect 5628 23102 5630 23154
rect 5682 23102 5908 23154
rect 5628 23100 5908 23102
rect 5628 23090 5684 23100
rect 5628 22932 5684 22942
rect 5628 21810 5684 22876
rect 5628 21758 5630 21810
rect 5682 21758 5684 21810
rect 5628 21746 5684 21758
rect 5852 21810 5908 23100
rect 6076 22372 6132 24668
rect 6412 24052 6468 25788
rect 7084 25732 7140 26796
rect 7420 26068 7476 26078
rect 7084 25730 7364 25732
rect 7084 25678 7086 25730
rect 7138 25678 7364 25730
rect 7084 25676 7364 25678
rect 7084 25666 7140 25676
rect 6860 25396 6916 25406
rect 6860 25302 6916 25340
rect 7308 24948 7364 25676
rect 7420 25730 7476 26012
rect 7420 25678 7422 25730
rect 7474 25678 7476 25730
rect 7420 25666 7476 25678
rect 7420 24948 7476 24958
rect 7308 24946 7476 24948
rect 7308 24894 7422 24946
rect 7474 24894 7476 24946
rect 7308 24892 7476 24894
rect 6636 24612 6692 24622
rect 6636 24518 6692 24556
rect 6076 22278 6132 22316
rect 6188 24050 6468 24052
rect 6188 23998 6414 24050
rect 6466 23998 6468 24050
rect 6188 23996 6468 23998
rect 5852 21758 5854 21810
rect 5906 21758 5908 21810
rect 5852 21746 5908 21758
rect 5292 20130 5684 20132
rect 5292 20078 5294 20130
rect 5346 20078 5684 20130
rect 5292 20076 5684 20078
rect 4956 19906 5012 19918
rect 4956 19854 4958 19906
rect 5010 19854 5012 19906
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4396 17892 4452 17902
rect 4396 17778 4452 17836
rect 4396 17726 4398 17778
rect 4450 17726 4452 17778
rect 4396 17714 4452 17726
rect 1708 17556 1764 17566
rect 1708 17462 1764 17500
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4956 16436 5012 19854
rect 5180 18564 5236 18574
rect 5292 18564 5348 20076
rect 5628 19234 5684 20076
rect 5852 20020 5908 20030
rect 5852 19926 5908 19964
rect 5628 19182 5630 19234
rect 5682 19182 5684 19234
rect 5628 19170 5684 19182
rect 5964 19010 6020 19022
rect 5964 18958 5966 19010
rect 6018 18958 6020 19010
rect 5964 18676 6020 18958
rect 5964 18610 6020 18620
rect 5180 18562 5348 18564
rect 5180 18510 5182 18562
rect 5234 18510 5348 18562
rect 5180 18508 5348 18510
rect 5180 18498 5236 18508
rect 6076 18452 6132 18462
rect 6076 18358 6132 18396
rect 5068 18226 5124 18238
rect 5068 18174 5070 18226
rect 5122 18174 5124 18226
rect 5068 17668 5124 18174
rect 5068 17574 5124 17612
rect 5740 17668 5796 17678
rect 5740 17574 5796 17612
rect 6076 17220 6132 17230
rect 5180 17108 5236 17118
rect 5516 17108 5572 17118
rect 5180 17106 5516 17108
rect 5180 17054 5182 17106
rect 5234 17054 5516 17106
rect 5180 17052 5516 17054
rect 5180 17042 5236 17052
rect 5516 17014 5572 17052
rect 6076 17106 6132 17164
rect 6076 17054 6078 17106
rect 6130 17054 6132 17106
rect 6076 17042 6132 17054
rect 6188 16770 6244 23996
rect 6412 23986 6468 23996
rect 7308 23940 7364 23950
rect 6524 23042 6580 23054
rect 6524 22990 6526 23042
rect 6578 22990 6580 23042
rect 6524 21924 6580 22990
rect 7196 23042 7252 23054
rect 7196 22990 7198 23042
rect 7250 22990 7252 23042
rect 7196 22932 7252 22990
rect 7196 22866 7252 22876
rect 6524 21858 6580 21868
rect 6636 22370 6692 22382
rect 6636 22318 6638 22370
rect 6690 22318 6692 22370
rect 6524 21700 6580 21710
rect 6412 21644 6524 21700
rect 6412 21586 6468 21644
rect 6412 21534 6414 21586
rect 6466 21534 6468 21586
rect 6412 21522 6468 21534
rect 6300 20692 6356 20702
rect 6300 20598 6356 20636
rect 6524 19234 6580 21644
rect 6636 21588 6692 22318
rect 6972 22372 7028 22382
rect 6972 22278 7028 22316
rect 6636 21522 6692 21532
rect 6748 22148 6804 22158
rect 6748 20132 6804 22092
rect 7308 21812 7364 23884
rect 7420 22372 7476 24892
rect 7532 22484 7588 27020
rect 8092 26290 8148 27132
rect 8092 26238 8094 26290
rect 8146 26238 8148 26290
rect 8092 25508 8148 26238
rect 8092 25442 8148 25452
rect 8204 27074 8260 27580
rect 8316 27570 8372 27580
rect 8876 27580 9044 27636
rect 8540 27300 8596 27310
rect 8540 27186 8596 27244
rect 8540 27134 8542 27186
rect 8594 27134 8596 27186
rect 8540 27122 8596 27134
rect 8204 27022 8206 27074
rect 8258 27022 8260 27074
rect 7868 24724 7924 24734
rect 7868 24612 7924 24668
rect 7756 24610 7924 24612
rect 7756 24558 7870 24610
rect 7922 24558 7924 24610
rect 7756 24556 7924 24558
rect 7756 23266 7812 24556
rect 7868 24546 7924 24556
rect 8204 23940 8260 27022
rect 8652 26178 8708 26190
rect 8652 26126 8654 26178
rect 8706 26126 8708 26178
rect 8652 25508 8708 26126
rect 8652 25442 8708 25452
rect 8540 24724 8596 24734
rect 8540 24630 8596 24668
rect 8204 23874 8260 23884
rect 8428 23938 8484 23950
rect 8428 23886 8430 23938
rect 8482 23886 8484 23938
rect 7756 23214 7758 23266
rect 7810 23214 7812 23266
rect 7756 23202 7812 23214
rect 8428 23154 8484 23886
rect 8428 23102 8430 23154
rect 8482 23102 8484 23154
rect 7756 23042 7812 23054
rect 7756 22990 7758 23042
rect 7810 22990 7812 23042
rect 7532 22428 7700 22484
rect 7420 22306 7476 22316
rect 7532 22258 7588 22270
rect 7532 22206 7534 22258
rect 7586 22206 7588 22258
rect 7532 22148 7588 22206
rect 7532 22082 7588 22092
rect 7196 21756 7364 21812
rect 6972 21474 7028 21486
rect 6972 21422 6974 21474
rect 7026 21422 7028 21474
rect 6972 20914 7028 21422
rect 6972 20862 6974 20914
rect 7026 20862 7028 20914
rect 6972 20244 7028 20862
rect 6972 20178 7028 20188
rect 6524 19182 6526 19234
rect 6578 19182 6580 19234
rect 6524 18564 6580 19182
rect 6524 18498 6580 18508
rect 6636 20076 6804 20132
rect 6524 18340 6580 18350
rect 6636 18340 6692 20076
rect 7084 20020 7140 20030
rect 6748 19964 7084 20020
rect 6748 19458 6804 19964
rect 7084 19926 7140 19964
rect 6748 19406 6750 19458
rect 6802 19406 6804 19458
rect 6748 19394 6804 19406
rect 7084 19348 7140 19358
rect 6860 19292 7084 19348
rect 6524 18338 6692 18340
rect 6524 18286 6526 18338
rect 6578 18286 6692 18338
rect 6524 18284 6692 18286
rect 6748 19236 6804 19246
rect 6748 18452 6804 19180
rect 6524 18274 6580 18284
rect 6524 17556 6580 17566
rect 6524 17554 6692 17556
rect 6524 17502 6526 17554
rect 6578 17502 6692 17554
rect 6524 17500 6692 17502
rect 6524 17490 6580 17500
rect 6188 16718 6190 16770
rect 6242 16718 6244 16770
rect 6188 16706 6244 16718
rect 6524 16770 6580 16782
rect 6524 16718 6526 16770
rect 6578 16718 6580 16770
rect 4284 16322 4340 16334
rect 4284 16270 4286 16322
rect 4338 16270 4340 16322
rect 4284 16210 4340 16270
rect 4956 16322 5012 16380
rect 4956 16270 4958 16322
rect 5010 16270 5012 16322
rect 4956 16258 5012 16270
rect 5180 16658 5236 16670
rect 5180 16606 5182 16658
rect 5234 16606 5236 16658
rect 4284 16158 4286 16210
rect 4338 16158 4340 16210
rect 4284 16146 4340 16158
rect 5180 16210 5236 16606
rect 5180 16158 5182 16210
rect 5234 16158 5236 16210
rect 4732 15988 4788 15998
rect 4732 15894 4788 15932
rect 5068 15540 5124 15550
rect 5068 15446 5124 15484
rect 5180 15148 5236 16158
rect 5516 16436 5572 16446
rect 5516 15538 5572 16380
rect 5516 15486 5518 15538
rect 5570 15486 5572 15538
rect 5516 15474 5572 15486
rect 5852 15986 5908 15998
rect 5852 15934 5854 15986
rect 5906 15934 5908 15986
rect 5180 15092 5460 15148
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 5180 14644 5236 14654
rect 5180 14550 5236 14588
rect 5404 14420 5460 15092
rect 5852 14868 5908 15934
rect 5964 15652 6020 15662
rect 5964 15538 6020 15596
rect 5964 15486 5966 15538
rect 6018 15486 6020 15538
rect 5964 15474 6020 15486
rect 5852 14644 5908 14812
rect 6412 15202 6468 15214
rect 6412 15150 6414 15202
rect 6466 15150 6468 15202
rect 6412 14756 6468 15150
rect 6524 15148 6580 16718
rect 6636 16324 6692 17500
rect 6748 16884 6804 18396
rect 6860 18450 6916 19292
rect 7084 19282 7140 19292
rect 6860 18398 6862 18450
rect 6914 18398 6916 18450
rect 6860 18004 6916 18398
rect 6860 16996 6916 17948
rect 7084 19124 7140 19134
rect 6972 17332 7028 17342
rect 6972 17106 7028 17276
rect 6972 17054 6974 17106
rect 7026 17054 7028 17106
rect 6972 17042 7028 17054
rect 7084 17108 7140 19068
rect 7196 18562 7252 21756
rect 7308 21588 7364 21598
rect 7308 21494 7364 21532
rect 7532 20802 7588 20814
rect 7532 20750 7534 20802
rect 7586 20750 7588 20802
rect 7308 20132 7364 20142
rect 7308 19236 7364 20076
rect 7532 20020 7588 20750
rect 7308 19170 7364 19180
rect 7420 19906 7476 19918
rect 7420 19854 7422 19906
rect 7474 19854 7476 19906
rect 7308 18676 7364 18686
rect 7420 18676 7476 19854
rect 7532 19236 7588 19964
rect 7644 19906 7700 22428
rect 7644 19854 7646 19906
rect 7698 19854 7700 19906
rect 7644 19842 7700 19854
rect 7756 19348 7812 22990
rect 8092 22148 8148 22158
rect 8316 22148 8372 22158
rect 7868 22146 8148 22148
rect 7868 22094 8094 22146
rect 8146 22094 8148 22146
rect 7868 22092 8148 22094
rect 7868 21476 7924 22092
rect 8092 22082 8148 22092
rect 8204 22146 8372 22148
rect 8204 22094 8318 22146
rect 8370 22094 8372 22146
rect 8204 22092 8372 22094
rect 8092 21588 8148 21598
rect 7868 21410 7924 21420
rect 7980 21474 8036 21486
rect 7980 21422 7982 21474
rect 8034 21422 8036 21474
rect 7980 20244 8036 21422
rect 7980 20178 8036 20188
rect 8092 20802 8148 21532
rect 8092 20750 8094 20802
rect 8146 20750 8148 20802
rect 8092 20020 8148 20750
rect 7756 19282 7812 19292
rect 7868 19964 8092 20020
rect 7644 19236 7700 19246
rect 7532 19234 7700 19236
rect 7532 19182 7646 19234
rect 7698 19182 7700 19234
rect 7532 19180 7700 19182
rect 7644 19170 7700 19180
rect 7868 19234 7924 19964
rect 8092 19954 8148 19964
rect 7868 19182 7870 19234
rect 7922 19182 7924 19234
rect 7868 19170 7924 19182
rect 7756 19012 7812 19022
rect 7308 18674 7476 18676
rect 7308 18622 7310 18674
rect 7362 18622 7476 18674
rect 7308 18620 7476 18622
rect 7308 18610 7364 18620
rect 7196 18510 7198 18562
rect 7250 18510 7252 18562
rect 7196 17666 7252 18510
rect 7196 17614 7198 17666
rect 7250 17614 7252 17666
rect 7196 17602 7252 17614
rect 7308 17668 7364 17678
rect 7084 17042 7140 17052
rect 6860 16930 6916 16940
rect 7196 16884 7252 16894
rect 7308 16884 7364 17612
rect 7420 17108 7476 18620
rect 7644 19010 7812 19012
rect 7644 18958 7758 19010
rect 7810 18958 7812 19010
rect 7644 18956 7812 18958
rect 7420 17042 7476 17052
rect 7532 18450 7588 18462
rect 7532 18398 7534 18450
rect 7586 18398 7588 18450
rect 6748 16818 6804 16828
rect 7084 16882 7364 16884
rect 7084 16830 7198 16882
rect 7250 16830 7364 16882
rect 7084 16828 7364 16830
rect 7084 16548 7140 16828
rect 7196 16818 7252 16828
rect 6636 16258 6692 16268
rect 6860 16492 7140 16548
rect 6524 15092 6804 15148
rect 5852 14578 5908 14588
rect 6076 14700 6468 14756
rect 6636 14980 6692 14990
rect 5404 14354 5460 14364
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 6076 13076 6132 14700
rect 6636 14642 6692 14924
rect 6636 14590 6638 14642
rect 6690 14590 6692 14642
rect 6636 14578 6692 14590
rect 6188 14532 6244 14542
rect 6188 13970 6244 14476
rect 6188 13918 6190 13970
rect 6242 13918 6244 13970
rect 6188 13906 6244 13918
rect 6524 14420 6580 14430
rect 6188 13076 6244 13086
rect 6076 13020 6188 13076
rect 6188 13010 6244 13020
rect 6524 13074 6580 14364
rect 6636 13748 6692 13758
rect 6636 13654 6692 13692
rect 6524 13022 6526 13074
rect 6578 13022 6580 13074
rect 6524 13010 6580 13022
rect 6748 12852 6804 15092
rect 6748 12786 6804 12796
rect 6860 13746 6916 16492
rect 7420 16436 7476 16446
rect 6972 16098 7028 16110
rect 6972 16046 6974 16098
rect 7026 16046 7028 16098
rect 6972 15764 7028 16046
rect 7420 16098 7476 16380
rect 7420 16046 7422 16098
rect 7474 16046 7476 16098
rect 7420 16034 7476 16046
rect 7532 16100 7588 18398
rect 7532 16006 7588 16044
rect 7644 16098 7700 18956
rect 7756 18946 7812 18956
rect 8204 18900 8260 22092
rect 8316 22082 8372 22092
rect 8428 21700 8484 23102
rect 8540 22372 8596 22382
rect 8540 22278 8596 22316
rect 8428 21634 8484 21644
rect 8876 20916 8932 27580
rect 8988 26964 9044 27002
rect 9212 26964 9268 28366
rect 9772 28642 9828 28654
rect 9772 28590 9774 28642
rect 9826 28590 9828 28642
rect 9548 27972 9604 27982
rect 9548 27878 9604 27916
rect 9772 27860 9828 28590
rect 10108 28644 10164 28654
rect 10108 28550 10164 28588
rect 9884 27972 9940 27982
rect 9884 27878 9940 27916
rect 9772 27794 9828 27804
rect 10444 27412 10500 29260
rect 11004 29204 11060 29214
rect 10556 28756 10612 28766
rect 10556 28642 10612 28700
rect 10556 28590 10558 28642
rect 10610 28590 10612 28642
rect 10556 28578 10612 28590
rect 10892 27972 10948 27982
rect 10444 27346 10500 27356
rect 10556 27858 10612 27870
rect 10780 27860 10836 27870
rect 10556 27806 10558 27858
rect 10610 27806 10612 27858
rect 9044 26908 9268 26964
rect 9548 27188 9604 27198
rect 8988 26898 9044 26908
rect 9436 26292 9492 26302
rect 9324 25732 9380 25770
rect 9324 25666 9380 25676
rect 9324 25508 9380 25518
rect 9324 25394 9380 25452
rect 9436 25506 9492 26236
rect 9436 25454 9438 25506
rect 9490 25454 9492 25506
rect 9436 25442 9492 25454
rect 9324 25342 9326 25394
rect 9378 25342 9380 25394
rect 9324 25330 9380 25342
rect 8988 25282 9044 25294
rect 8988 25230 8990 25282
rect 9042 25230 9044 25282
rect 8988 25172 9044 25230
rect 8988 25106 9044 25116
rect 9548 24948 9604 27132
rect 10444 27076 10500 27086
rect 10556 27076 10612 27806
rect 10500 27020 10612 27076
rect 10668 27804 10780 27860
rect 10668 27074 10724 27804
rect 10780 27766 10836 27804
rect 10668 27022 10670 27074
rect 10722 27022 10724 27074
rect 10444 26982 10500 27020
rect 10108 26292 10164 26302
rect 10332 26292 10388 26302
rect 10108 26198 10164 26236
rect 10220 26290 10388 26292
rect 10220 26238 10334 26290
rect 10386 26238 10388 26290
rect 10220 26236 10388 26238
rect 9772 26178 9828 26190
rect 9772 26126 9774 26178
rect 9826 26126 9828 26178
rect 9772 25284 9828 26126
rect 10220 25620 10276 26236
rect 10332 26226 10388 26236
rect 10668 26292 10724 27022
rect 10780 27076 10836 27086
rect 10892 27076 10948 27916
rect 11004 27858 11060 29148
rect 12460 29204 12516 30718
rect 13916 30436 13972 30446
rect 13692 30212 13748 30222
rect 13692 30118 13748 30156
rect 13916 30098 13972 30380
rect 15484 30436 15540 30942
rect 16156 30994 16212 31164
rect 16604 31154 16660 31164
rect 16716 32562 16772 32574
rect 16716 32510 16718 32562
rect 16770 32510 16772 32562
rect 16716 31108 16772 32510
rect 18508 31666 18564 32620
rect 18508 31614 18510 31666
rect 18562 31614 18564 31666
rect 18508 31602 18564 31614
rect 17500 31556 17556 31566
rect 17500 31218 17556 31500
rect 18172 31556 18228 31566
rect 18956 31556 19012 31566
rect 19068 31556 19124 33070
rect 18228 31500 18452 31556
rect 18172 31462 18228 31500
rect 17500 31166 17502 31218
rect 17554 31166 17556 31218
rect 17500 31154 17556 31166
rect 17836 31220 17892 31230
rect 16716 31042 16772 31052
rect 17836 31106 17892 31164
rect 17836 31054 17838 31106
rect 17890 31054 17892 31106
rect 17836 30996 17892 31054
rect 16156 30942 16158 30994
rect 16210 30942 16212 30994
rect 16156 30930 16212 30942
rect 17500 30940 17892 30996
rect 15484 30370 15540 30380
rect 17052 30548 17108 30558
rect 13916 30046 13918 30098
rect 13970 30046 13972 30098
rect 13916 30034 13972 30046
rect 16940 30100 16996 30110
rect 16940 30006 16996 30044
rect 13916 29708 14196 29764
rect 13692 29652 13748 29662
rect 13916 29652 13972 29708
rect 13692 29650 13972 29652
rect 13692 29598 13694 29650
rect 13746 29598 13972 29650
rect 13692 29596 13972 29598
rect 13692 29586 13748 29596
rect 12460 29138 12516 29148
rect 14028 29538 14084 29550
rect 14028 29486 14030 29538
rect 14082 29486 14084 29538
rect 12012 28868 12068 28878
rect 12012 28642 12068 28812
rect 12012 28590 12014 28642
rect 12066 28590 12068 28642
rect 12012 28578 12068 28590
rect 13468 28868 13524 28878
rect 13468 28642 13524 28812
rect 13468 28590 13470 28642
rect 13522 28590 13524 28642
rect 13468 28578 13524 28590
rect 13580 28644 13636 28654
rect 13916 28644 13972 28654
rect 13580 28642 13916 28644
rect 13580 28590 13582 28642
rect 13634 28590 13916 28642
rect 13580 28588 13916 28590
rect 13580 28578 13636 28588
rect 11564 28532 11620 28542
rect 11452 28530 11620 28532
rect 11452 28478 11566 28530
rect 11618 28478 11620 28530
rect 11452 28476 11620 28478
rect 11004 27806 11006 27858
rect 11058 27806 11060 27858
rect 11004 27794 11060 27806
rect 11228 27972 11284 27982
rect 11228 27858 11284 27916
rect 11228 27806 11230 27858
rect 11282 27806 11284 27858
rect 11228 27794 11284 27806
rect 11228 27524 11284 27534
rect 10780 27074 10892 27076
rect 10780 27022 10782 27074
rect 10834 27022 10892 27074
rect 10780 27020 10892 27022
rect 10780 27010 10836 27020
rect 10892 26982 10948 27020
rect 11004 27412 11060 27422
rect 11004 26908 11060 27356
rect 10668 26226 10724 26236
rect 10780 26852 11060 26908
rect 11116 27300 11172 27310
rect 9884 25564 10276 25620
rect 10556 25732 10612 25742
rect 9884 25508 9940 25564
rect 9884 25414 9940 25452
rect 9884 25284 9940 25294
rect 9772 25228 9884 25284
rect 9436 24892 9604 24948
rect 8988 24836 9044 24846
rect 8988 24742 9044 24780
rect 9324 23940 9380 23950
rect 9436 23940 9492 24892
rect 9324 23938 9492 23940
rect 9324 23886 9326 23938
rect 9378 23886 9492 23938
rect 9324 23884 9492 23886
rect 9548 24724 9604 24734
rect 9548 23940 9604 24668
rect 9660 23940 9716 23950
rect 9548 23938 9716 23940
rect 9548 23886 9662 23938
rect 9714 23886 9716 23938
rect 9548 23884 9716 23886
rect 9324 23156 9380 23884
rect 9660 23874 9716 23884
rect 9324 23090 9380 23100
rect 9884 23044 9940 25228
rect 10108 24722 10164 25564
rect 10556 25508 10612 25676
rect 10668 25508 10724 25518
rect 10556 25506 10724 25508
rect 10556 25454 10670 25506
rect 10722 25454 10724 25506
rect 10556 25452 10724 25454
rect 10332 25396 10388 25406
rect 10332 25394 10500 25396
rect 10332 25342 10334 25394
rect 10386 25342 10500 25394
rect 10332 25340 10500 25342
rect 10332 25330 10388 25340
rect 10108 24670 10110 24722
rect 10162 24670 10164 24722
rect 10108 24658 10164 24670
rect 9996 23828 10052 23838
rect 9996 23734 10052 23772
rect 10220 23154 10276 23166
rect 10220 23102 10222 23154
rect 10274 23102 10276 23154
rect 9996 23044 10052 23054
rect 9884 23042 10052 23044
rect 9884 22990 9998 23042
rect 10050 22990 10052 23042
rect 9884 22988 10052 22990
rect 9884 22484 9940 22494
rect 8988 22372 9044 22382
rect 8988 22278 9044 22316
rect 9324 22146 9380 22158
rect 9324 22094 9326 22146
rect 9378 22094 9380 22146
rect 8988 21476 9044 21486
rect 9044 21420 9156 21476
rect 8988 21382 9044 21420
rect 8988 20916 9044 20926
rect 8876 20914 9044 20916
rect 8876 20862 8990 20914
rect 9042 20862 9044 20914
rect 8876 20860 9044 20862
rect 8316 20804 8372 20814
rect 8316 19234 8372 20748
rect 8652 20690 8708 20702
rect 8652 20638 8654 20690
rect 8706 20638 8708 20690
rect 8652 20580 8708 20638
rect 8540 20020 8596 20030
rect 8540 19926 8596 19964
rect 8316 19182 8318 19234
rect 8370 19182 8372 19234
rect 8316 19170 8372 19182
rect 8428 19906 8484 19918
rect 8428 19854 8430 19906
rect 8482 19854 8484 19906
rect 7868 18844 8260 18900
rect 7868 18450 7924 18844
rect 7980 18676 8036 18686
rect 7980 18562 8036 18620
rect 7980 18510 7982 18562
rect 8034 18510 8036 18562
rect 7980 18498 8036 18510
rect 8316 18564 8372 18574
rect 8316 18470 8372 18508
rect 7868 18398 7870 18450
rect 7922 18398 7924 18450
rect 7756 17780 7812 17790
rect 7756 17686 7812 17724
rect 7756 17108 7812 17118
rect 7756 17014 7812 17052
rect 7644 16046 7646 16098
rect 7698 16046 7700 16098
rect 7644 15764 7700 16046
rect 6972 15708 7700 15764
rect 7756 16884 7812 16894
rect 7756 15652 7812 16828
rect 7532 15596 7812 15652
rect 7084 15426 7140 15438
rect 7084 15374 7086 15426
rect 7138 15374 7140 15426
rect 7084 15148 7140 15374
rect 7308 15316 7364 15326
rect 7308 15148 7364 15260
rect 7084 15092 7364 15148
rect 7196 14644 7252 14654
rect 6972 14588 7196 14644
rect 6972 14530 7028 14588
rect 6972 14478 6974 14530
rect 7026 14478 7028 14530
rect 6972 14466 7028 14478
rect 6860 13694 6862 13746
rect 6914 13694 6916 13746
rect 6860 12516 6916 13694
rect 7084 13746 7140 14588
rect 7196 14578 7252 14588
rect 7308 14642 7364 15092
rect 7308 14590 7310 14642
rect 7362 14590 7364 14642
rect 7308 14578 7364 14590
rect 7420 14308 7476 14318
rect 7420 13970 7476 14252
rect 7420 13918 7422 13970
rect 7474 13918 7476 13970
rect 7420 13906 7476 13918
rect 7532 13748 7588 15596
rect 7644 15314 7700 15326
rect 7644 15262 7646 15314
rect 7698 15262 7700 15314
rect 7644 15204 7700 15262
rect 7644 15138 7700 15148
rect 7868 14644 7924 18398
rect 8092 17780 8148 17790
rect 8092 17108 8148 17724
rect 8428 17780 8484 19854
rect 8652 19012 8708 20524
rect 8764 19796 8820 19806
rect 8764 19702 8820 19740
rect 8988 19460 9044 20860
rect 9100 20468 9156 21420
rect 9324 20804 9380 22094
rect 9324 20738 9380 20748
rect 9772 21140 9828 21150
rect 9548 20578 9604 20590
rect 9548 20526 9550 20578
rect 9602 20526 9604 20578
rect 9212 20468 9268 20478
rect 9100 20412 9212 20468
rect 9268 20412 9380 20468
rect 9212 20402 9268 20412
rect 8988 19404 9268 19460
rect 9100 19236 9156 19246
rect 9100 19142 9156 19180
rect 8652 18946 8708 18956
rect 8988 19010 9044 19022
rect 9212 19012 9268 19404
rect 8988 18958 8990 19010
rect 9042 18958 9044 19010
rect 8988 18900 9044 18958
rect 8988 18834 9044 18844
rect 9100 18956 9268 19012
rect 8988 18676 9044 18686
rect 8876 18564 8932 18574
rect 8428 17714 8484 17724
rect 8652 17892 8708 17902
rect 8652 17778 8708 17836
rect 8652 17726 8654 17778
rect 8706 17726 8708 17778
rect 8652 17714 8708 17726
rect 8316 17668 8372 17678
rect 8316 17574 8372 17612
rect 8092 17106 8260 17108
rect 8092 17054 8094 17106
rect 8146 17054 8260 17106
rect 8092 17052 8260 17054
rect 8092 17042 8148 17052
rect 8092 15874 8148 15886
rect 8092 15822 8094 15874
rect 8146 15822 8148 15874
rect 8092 15764 8148 15822
rect 8092 15698 8148 15708
rect 8204 15540 8260 17052
rect 8652 16996 8708 17006
rect 8652 16902 8708 16940
rect 8876 16436 8932 18508
rect 8988 18562 9044 18620
rect 8988 18510 8990 18562
rect 9042 18510 9044 18562
rect 8988 18498 9044 18510
rect 8876 16380 9044 16436
rect 8876 16212 8932 16222
rect 8876 16098 8932 16156
rect 8876 16046 8878 16098
rect 8930 16046 8932 16098
rect 8876 16034 8932 16046
rect 7868 14530 7924 14588
rect 7868 14478 7870 14530
rect 7922 14478 7924 14530
rect 7868 14466 7924 14478
rect 8092 15484 8260 15540
rect 7756 13972 7812 13982
rect 7084 13694 7086 13746
rect 7138 13694 7140 13746
rect 7084 13682 7140 13694
rect 7420 13692 7588 13748
rect 7644 13916 7756 13972
rect 6972 12964 7028 12974
rect 6972 12870 7028 12908
rect 7308 12852 7364 12862
rect 7308 12758 7364 12796
rect 6860 12460 7364 12516
rect 7308 12404 7364 12460
rect 7308 12178 7364 12348
rect 7308 12126 7310 12178
rect 7362 12126 7364 12178
rect 7308 12114 7364 12126
rect 6636 12066 6692 12078
rect 6636 12014 6638 12066
rect 6690 12014 6692 12066
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 6636 11620 6692 12014
rect 6636 11554 6692 11564
rect 7084 12066 7140 12078
rect 7084 12014 7086 12066
rect 7138 12014 7140 12066
rect 7084 11508 7140 12014
rect 7084 11442 7140 11452
rect 7420 10836 7476 13692
rect 7532 12180 7588 12190
rect 7644 12180 7700 13916
rect 7756 13878 7812 13916
rect 7868 13412 7924 13422
rect 7868 13074 7924 13356
rect 7868 13022 7870 13074
rect 7922 13022 7924 13074
rect 7868 13010 7924 13022
rect 7532 12178 7700 12180
rect 7532 12126 7534 12178
rect 7586 12126 7700 12178
rect 7532 12124 7700 12126
rect 8092 12962 8148 15484
rect 8428 15426 8484 15438
rect 8428 15374 8430 15426
rect 8482 15374 8484 15426
rect 8428 15204 8484 15374
rect 8204 15148 8484 15204
rect 8764 15428 8820 15438
rect 8204 13636 8260 15148
rect 8316 14644 8372 14654
rect 8372 14588 8484 14644
rect 8316 14550 8372 14588
rect 8316 13972 8372 13982
rect 8316 13858 8372 13916
rect 8316 13806 8318 13858
rect 8370 13806 8372 13858
rect 8316 13794 8372 13806
rect 8204 13570 8260 13580
rect 8428 13524 8484 14588
rect 8652 14420 8708 14430
rect 8652 14326 8708 14364
rect 8764 13860 8820 15372
rect 8988 15316 9044 16380
rect 8876 15314 9044 15316
rect 8876 15262 8990 15314
rect 9042 15262 9044 15314
rect 8876 15260 9044 15262
rect 8876 13972 8932 15260
rect 8988 15250 9044 15260
rect 9100 15148 9156 18956
rect 9324 18676 9380 20412
rect 9548 20020 9604 20526
rect 9772 20130 9828 21084
rect 9772 20078 9774 20130
rect 9826 20078 9828 20130
rect 9772 20066 9828 20078
rect 9212 18620 9380 18676
rect 9436 20018 9604 20020
rect 9436 19966 9550 20018
rect 9602 19966 9604 20018
rect 9436 19964 9604 19966
rect 9436 18676 9492 19964
rect 9548 19954 9604 19964
rect 9660 19236 9716 19274
rect 9660 19170 9716 19180
rect 9884 19124 9940 22428
rect 9548 19012 9604 19022
rect 9548 18918 9604 18956
rect 9772 19010 9828 19022
rect 9772 18958 9774 19010
rect 9826 18958 9828 19010
rect 9212 18452 9268 18620
rect 9436 18610 9492 18620
rect 9772 18564 9828 18958
rect 9772 18498 9828 18508
rect 9212 18396 9380 18452
rect 8876 13878 8932 13916
rect 8988 15092 9156 15148
rect 9212 15988 9268 15998
rect 8092 12910 8094 12962
rect 8146 12910 8148 12962
rect 7532 11732 7588 12124
rect 7868 11956 7924 11966
rect 7868 11862 7924 11900
rect 7532 11666 7588 11676
rect 7756 11620 7812 11630
rect 7644 11564 7756 11620
rect 7532 11508 7588 11518
rect 7644 11508 7700 11564
rect 7756 11554 7812 11564
rect 7532 11506 7700 11508
rect 7532 11454 7534 11506
rect 7586 11454 7700 11506
rect 7532 11452 7700 11454
rect 7532 11442 7588 11452
rect 8092 11396 8148 12910
rect 8316 13468 8484 13524
rect 8652 13858 8820 13860
rect 8652 13806 8766 13858
rect 8818 13806 8820 13858
rect 8652 13804 8820 13806
rect 8204 12404 8260 12414
rect 8204 12310 8260 12348
rect 8316 11956 8372 13468
rect 8652 13076 8708 13804
rect 8764 13794 8820 13804
rect 8988 13188 9044 15092
rect 9100 13972 9156 13982
rect 9100 13878 9156 13916
rect 8988 13132 9156 13188
rect 8652 13074 9044 13076
rect 8652 13022 8654 13074
rect 8706 13022 9044 13074
rect 8652 13020 9044 13022
rect 8652 13010 8708 13020
rect 8988 12962 9044 13020
rect 8988 12910 8990 12962
rect 9042 12910 9044 12962
rect 8988 12898 9044 12910
rect 8092 11330 8148 11340
rect 8204 11900 8372 11956
rect 8652 12852 8708 12862
rect 8092 11172 8148 11182
rect 8204 11172 8260 11900
rect 8316 11732 8372 11742
rect 8372 11676 8484 11732
rect 8316 11666 8372 11676
rect 8428 11394 8484 11676
rect 8428 11342 8430 11394
rect 8482 11342 8484 11394
rect 8428 11330 8484 11342
rect 8092 11170 8260 11172
rect 8092 11118 8094 11170
rect 8146 11118 8260 11170
rect 8092 11116 8260 11118
rect 8092 11106 8148 11116
rect 7420 10770 7476 10780
rect 8204 10836 8260 10846
rect 8204 10742 8260 10780
rect 8652 10834 8708 12796
rect 8764 12180 8820 12190
rect 8764 12086 8820 12124
rect 9100 11732 9156 13132
rect 8652 10782 8654 10834
rect 8706 10782 8708 10834
rect 8652 10770 8708 10782
rect 8764 11676 9156 11732
rect 8764 11060 8820 11676
rect 9212 11620 9268 15932
rect 9324 14308 9380 18396
rect 9772 18340 9828 18378
rect 9772 18274 9828 18284
rect 9772 18116 9828 18126
rect 9772 17890 9828 18060
rect 9772 17838 9774 17890
rect 9826 17838 9828 17890
rect 9772 17826 9828 17838
rect 9772 17332 9828 17342
rect 9660 16324 9716 16334
rect 9548 16100 9604 16110
rect 9548 15538 9604 16044
rect 9548 15486 9550 15538
rect 9602 15486 9604 15538
rect 9548 15474 9604 15486
rect 9324 14242 9380 14252
rect 9660 14530 9716 16268
rect 9660 14478 9662 14530
rect 9714 14478 9716 14530
rect 9660 12404 9716 14478
rect 9660 12338 9716 12348
rect 9772 16210 9828 17276
rect 9772 16158 9774 16210
rect 9826 16158 9828 16210
rect 9772 11620 9828 16158
rect 9884 16100 9940 19068
rect 9996 17556 10052 22988
rect 10108 22932 10164 22942
rect 10220 22932 10276 23102
rect 10164 22876 10276 22932
rect 10108 22484 10164 22876
rect 10108 22482 10388 22484
rect 10108 22430 10110 22482
rect 10162 22430 10388 22482
rect 10108 22428 10388 22430
rect 10108 22418 10164 22428
rect 10332 21810 10388 22428
rect 10332 21758 10334 21810
rect 10386 21758 10388 21810
rect 10332 21746 10388 21758
rect 10108 21474 10164 21486
rect 10108 21422 10110 21474
rect 10162 21422 10164 21474
rect 10108 20692 10164 21422
rect 10220 20804 10276 20814
rect 10220 20710 10276 20748
rect 10108 18340 10164 20636
rect 10108 18274 10164 18284
rect 10220 19906 10276 19918
rect 10220 19854 10222 19906
rect 10274 19854 10276 19906
rect 10220 19348 10276 19854
rect 9996 17490 10052 17500
rect 10108 17668 10164 17678
rect 10108 17106 10164 17612
rect 10108 17054 10110 17106
rect 10162 17054 10164 17106
rect 10108 17042 10164 17054
rect 9884 16034 9940 16044
rect 9996 16884 10052 16894
rect 9996 15202 10052 16828
rect 10220 15204 10276 19292
rect 10444 18900 10500 25340
rect 10556 22370 10612 25452
rect 10668 25442 10724 25452
rect 10780 23156 10836 26852
rect 11004 25508 11060 25518
rect 11004 25414 11060 25452
rect 11004 24610 11060 24622
rect 11004 24558 11006 24610
rect 11058 24558 11060 24610
rect 11004 24500 11060 24558
rect 11004 24434 11060 24444
rect 11004 23938 11060 23950
rect 11004 23886 11006 23938
rect 11058 23886 11060 23938
rect 11004 23380 11060 23886
rect 11004 23314 11060 23324
rect 10556 22318 10558 22370
rect 10610 22318 10612 22370
rect 10556 22306 10612 22318
rect 10668 23100 10836 23156
rect 11004 23156 11060 23166
rect 10668 19460 10724 23100
rect 11004 23062 11060 23100
rect 10892 23044 10948 23054
rect 10780 23042 10948 23044
rect 10780 22990 10894 23042
rect 10946 22990 10948 23042
rect 10780 22988 10948 22990
rect 10780 20804 10836 22988
rect 10892 22978 10948 22988
rect 10892 21476 10948 21486
rect 10892 21382 10948 21420
rect 10780 20738 10836 20748
rect 11116 20468 11172 27244
rect 11228 27298 11284 27468
rect 11228 27246 11230 27298
rect 11282 27246 11284 27298
rect 11228 27234 11284 27246
rect 11452 26908 11508 28476
rect 11564 28466 11620 28476
rect 13020 28418 13076 28430
rect 13020 28366 13022 28418
rect 13074 28366 13076 28418
rect 12348 27972 12404 27982
rect 12348 27858 12404 27916
rect 12348 27806 12350 27858
rect 12402 27806 12404 27858
rect 12348 27794 12404 27806
rect 12124 27748 12180 27758
rect 12124 27746 12292 27748
rect 12124 27694 12126 27746
rect 12178 27694 12292 27746
rect 12124 27692 12292 27694
rect 12124 27682 12180 27692
rect 11676 27636 11732 27646
rect 11676 27542 11732 27580
rect 12236 27188 12292 27692
rect 11564 27076 11620 27114
rect 11564 27010 11620 27020
rect 12124 26964 12180 27002
rect 11452 26852 11620 26908
rect 12124 26898 12180 26908
rect 11340 25730 11396 25742
rect 11340 25678 11342 25730
rect 11394 25678 11396 25730
rect 11340 25396 11396 25678
rect 11340 25330 11396 25340
rect 11452 25508 11508 25518
rect 11452 24836 11508 25452
rect 11340 23826 11396 23838
rect 11340 23774 11342 23826
rect 11394 23774 11396 23826
rect 11340 23268 11396 23774
rect 11340 22036 11396 23212
rect 11340 21970 11396 21980
rect 11452 22820 11508 24780
rect 11564 22932 11620 26852
rect 12236 26290 12292 27132
rect 12684 27634 12740 27646
rect 12684 27582 12686 27634
rect 12738 27582 12740 27634
rect 12684 27076 12740 27582
rect 12908 27076 12964 27086
rect 12684 27020 12908 27076
rect 12908 26982 12964 27020
rect 12236 26238 12238 26290
rect 12290 26238 12292 26290
rect 12236 26226 12292 26238
rect 12460 26740 12516 26750
rect 11676 26178 11732 26190
rect 11676 26126 11678 26178
rect 11730 26126 11732 26178
rect 11676 25620 11732 26126
rect 12124 25956 12180 25966
rect 11676 25554 11732 25564
rect 11900 25732 11956 25742
rect 11900 25618 11956 25676
rect 11900 25566 11902 25618
rect 11954 25566 11956 25618
rect 11900 25554 11956 25566
rect 11788 25396 11844 25406
rect 11788 23828 11844 25340
rect 12012 25284 12068 25294
rect 11900 24948 11956 24958
rect 11900 24612 11956 24892
rect 12012 24834 12068 25228
rect 12012 24782 12014 24834
rect 12066 24782 12068 24834
rect 12012 24770 12068 24782
rect 11900 23938 11956 24556
rect 11900 23886 11902 23938
rect 11954 23886 11956 23938
rect 11900 23874 11956 23886
rect 11564 22866 11620 22876
rect 11676 23380 11732 23390
rect 11676 23266 11732 23324
rect 11676 23214 11678 23266
rect 11730 23214 11732 23266
rect 11228 21812 11284 21822
rect 11452 21812 11508 22764
rect 11676 22372 11732 23214
rect 11676 22306 11732 22316
rect 11564 22258 11620 22270
rect 11564 22206 11566 22258
rect 11618 22206 11620 22258
rect 11564 21924 11620 22206
rect 11564 21858 11620 21868
rect 11676 22036 11732 22046
rect 11228 21586 11284 21756
rect 11228 21534 11230 21586
rect 11282 21534 11284 21586
rect 11228 21522 11284 21534
rect 11340 21756 11508 21812
rect 11340 21364 11396 21756
rect 11564 21700 11620 21710
rect 10668 19394 10724 19404
rect 10780 20412 11172 20468
rect 11228 21308 11396 21364
rect 11452 21644 11564 21700
rect 10444 18844 10724 18900
rect 10556 18676 10612 18686
rect 10332 18564 10388 18574
rect 10332 18470 10388 18508
rect 10444 18452 10500 18490
rect 10444 18386 10500 18396
rect 10444 18228 10500 18238
rect 10332 18004 10388 18014
rect 10332 16996 10388 17948
rect 10332 16210 10388 16940
rect 10332 16158 10334 16210
rect 10386 16158 10388 16210
rect 10332 16146 10388 16158
rect 10444 16098 10500 18172
rect 10556 17106 10612 18620
rect 10668 17778 10724 18844
rect 10668 17726 10670 17778
rect 10722 17726 10724 17778
rect 10668 17714 10724 17726
rect 10780 17666 10836 20412
rect 10892 20018 10948 20030
rect 10892 19966 10894 20018
rect 10946 19966 10948 20018
rect 10892 19684 10948 19966
rect 10892 19628 11172 19684
rect 11004 19460 11060 19470
rect 10780 17614 10782 17666
rect 10834 17614 10836 17666
rect 10556 17054 10558 17106
rect 10610 17054 10612 17106
rect 10556 17042 10612 17054
rect 10668 17556 10724 17566
rect 10444 16046 10446 16098
rect 10498 16046 10500 16098
rect 10444 15988 10500 16046
rect 10444 15922 10500 15932
rect 9996 15150 9998 15202
rect 10050 15150 10052 15202
rect 9996 15138 10052 15150
rect 10108 15148 10276 15204
rect 10668 15148 10724 17500
rect 10780 16882 10836 17614
rect 10780 16830 10782 16882
rect 10834 16830 10836 16882
rect 10780 16818 10836 16830
rect 10892 19124 10948 19134
rect 10780 16322 10836 16334
rect 10780 16270 10782 16322
rect 10834 16270 10836 16322
rect 10780 15538 10836 16270
rect 10780 15486 10782 15538
rect 10834 15486 10836 15538
rect 10780 15428 10836 15486
rect 10780 15362 10836 15372
rect 10108 13524 10164 15148
rect 10444 15092 10724 15148
rect 10220 13748 10276 13786
rect 10220 13682 10276 13692
rect 10332 13636 10388 13646
rect 10332 13542 10388 13580
rect 9996 13468 10164 13524
rect 10220 13524 10276 13534
rect 9996 12402 10052 13468
rect 9996 12350 9998 12402
rect 10050 12350 10052 12402
rect 9996 12338 10052 12350
rect 10108 13076 10164 13086
rect 9100 11564 9268 11620
rect 9660 11564 9828 11620
rect 8876 11284 8932 11294
rect 9100 11284 9156 11564
rect 9212 11396 9268 11406
rect 9212 11302 9268 11340
rect 8876 11282 9156 11284
rect 8876 11230 8878 11282
rect 8930 11230 9156 11282
rect 8876 11228 9156 11230
rect 8876 11218 8932 11228
rect 8764 10612 8820 11004
rect 8540 10556 8820 10612
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 8540 9938 8596 10556
rect 8540 9886 8542 9938
rect 8594 9886 8596 9938
rect 8540 9874 8596 9886
rect 8988 9716 9044 11228
rect 9100 10724 9156 10734
rect 9100 10630 9156 10668
rect 9436 9940 9492 9950
rect 9436 9846 9492 9884
rect 8988 9622 9044 9660
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 9660 7700 9716 11564
rect 9772 11396 9828 11406
rect 9772 9826 9828 11340
rect 10108 11172 10164 13020
rect 10220 12292 10276 13468
rect 10220 12198 10276 12236
rect 10444 11954 10500 15092
rect 10892 14980 10948 19068
rect 11004 18676 11060 19404
rect 11004 18610 11060 18620
rect 11116 18452 11172 19628
rect 11004 18396 11172 18452
rect 11004 18228 11060 18396
rect 11004 18162 11060 18172
rect 10668 14924 10948 14980
rect 11004 17778 11060 17790
rect 11004 17726 11006 17778
rect 11058 17726 11060 17778
rect 11004 17332 11060 17726
rect 11228 17554 11284 21308
rect 11340 20916 11396 20926
rect 11452 20916 11508 21644
rect 11564 21606 11620 21644
rect 11340 20914 11508 20916
rect 11340 20862 11342 20914
rect 11394 20862 11508 20914
rect 11340 20860 11508 20862
rect 11340 20850 11396 20860
rect 11564 20132 11620 20142
rect 11452 20020 11508 20030
rect 11340 19908 11396 19918
rect 11340 19814 11396 19852
rect 11452 19234 11508 19964
rect 11452 19182 11454 19234
rect 11506 19182 11508 19234
rect 11452 19170 11508 19182
rect 11564 19346 11620 20076
rect 11564 19294 11566 19346
rect 11618 19294 11620 19346
rect 11340 18676 11396 18686
rect 11340 18582 11396 18620
rect 11452 18564 11508 18574
rect 11340 18228 11396 18238
rect 11340 17780 11396 18172
rect 11340 17666 11396 17724
rect 11340 17614 11342 17666
rect 11394 17614 11396 17666
rect 11340 17602 11396 17614
rect 11228 17502 11230 17554
rect 11282 17502 11284 17554
rect 11228 17490 11284 17502
rect 11004 17276 11396 17332
rect 10556 14756 10612 14766
rect 10556 13858 10612 14700
rect 10556 13806 10558 13858
rect 10610 13806 10612 13858
rect 10556 13794 10612 13806
rect 10444 11902 10446 11954
rect 10498 11902 10500 11954
rect 10444 11732 10500 11902
rect 10668 11788 10724 14924
rect 11004 14530 11060 17276
rect 11004 14478 11006 14530
rect 11058 14478 11060 14530
rect 10892 14420 10948 14430
rect 10892 14326 10948 14364
rect 11004 13860 11060 14478
rect 10892 13804 11060 13860
rect 11116 17108 11172 17118
rect 10892 13524 10948 13804
rect 11004 13636 11060 13646
rect 11004 13542 11060 13580
rect 10892 13458 10948 13468
rect 11116 13412 11172 17052
rect 11340 16882 11396 17276
rect 11340 16830 11342 16882
rect 11394 16830 11396 16882
rect 11340 16818 11396 16830
rect 11228 16660 11284 16670
rect 11228 15538 11284 16604
rect 11228 15486 11230 15538
rect 11282 15486 11284 15538
rect 11228 15474 11284 15486
rect 11452 15540 11508 18508
rect 11564 17108 11620 19294
rect 11676 18900 11732 21980
rect 11788 21252 11844 23772
rect 12012 22258 12068 22270
rect 12012 22206 12014 22258
rect 12066 22206 12068 22258
rect 11788 21186 11844 21196
rect 11900 21474 11956 21486
rect 11900 21422 11902 21474
rect 11954 21422 11956 21474
rect 11788 20804 11844 20814
rect 11788 20710 11844 20748
rect 11900 20356 11956 21422
rect 12012 21028 12068 22206
rect 12012 20962 12068 20972
rect 11900 20290 11956 20300
rect 12012 20132 12068 20142
rect 12012 19236 12068 20076
rect 12012 19142 12068 19180
rect 12124 19012 12180 25900
rect 12236 25508 12292 25518
rect 12236 25414 12292 25452
rect 12460 25396 12516 26684
rect 12460 25302 12516 25340
rect 12684 26178 12740 26190
rect 12684 26126 12686 26178
rect 12738 26126 12740 26178
rect 12684 25508 12740 26126
rect 13020 26180 13076 28366
rect 13244 27970 13300 27982
rect 13244 27918 13246 27970
rect 13298 27918 13300 27970
rect 13244 27300 13300 27918
rect 13804 27970 13860 28588
rect 13916 28550 13972 28588
rect 14028 28196 14084 29486
rect 13804 27918 13806 27970
rect 13858 27918 13860 27970
rect 13804 27906 13860 27918
rect 13916 28140 14084 28196
rect 13244 27234 13300 27244
rect 13804 27300 13860 27310
rect 13020 26114 13076 26124
rect 13356 26964 13412 26974
rect 12684 24836 12740 25452
rect 12908 25394 12964 25406
rect 12908 25342 12910 25394
rect 12962 25342 12964 25394
rect 12908 24948 12964 25342
rect 13020 25396 13076 25406
rect 13020 25302 13076 25340
rect 12908 24882 12964 24892
rect 13020 24836 13076 24846
rect 12684 24834 12852 24836
rect 12684 24782 12686 24834
rect 12738 24782 12852 24834
rect 12684 24780 12852 24782
rect 12684 24770 12740 24780
rect 12684 24500 12740 24510
rect 12236 23042 12292 23054
rect 12236 22990 12238 23042
rect 12290 22990 12292 23042
rect 12236 22484 12292 22990
rect 12236 22418 12292 22428
rect 12460 22372 12516 22382
rect 12460 22278 12516 22316
rect 12348 21924 12404 21934
rect 12348 21252 12404 21868
rect 12460 21476 12516 21486
rect 12460 21474 12628 21476
rect 12460 21422 12462 21474
rect 12514 21422 12628 21474
rect 12460 21420 12628 21422
rect 12460 21410 12516 21420
rect 12572 21252 12628 21420
rect 12348 21196 12516 21252
rect 12236 21140 12292 21150
rect 12292 21084 12404 21140
rect 12236 21074 12292 21084
rect 12236 20914 12292 20926
rect 12236 20862 12238 20914
rect 12290 20862 12292 20914
rect 12236 20692 12292 20862
rect 12236 19124 12292 20636
rect 12236 19058 12292 19068
rect 11676 18834 11732 18844
rect 12012 18956 12180 19012
rect 11564 17042 11620 17052
rect 11676 17780 11732 17790
rect 11676 16770 11732 17724
rect 11676 16718 11678 16770
rect 11730 16718 11732 16770
rect 11676 16706 11732 16718
rect 11452 15426 11508 15484
rect 11452 15374 11454 15426
rect 11506 15374 11508 15426
rect 11452 15362 11508 15374
rect 11788 15540 11844 15550
rect 11788 15314 11844 15484
rect 12012 15426 12068 18956
rect 12348 16436 12404 21084
rect 12348 16098 12404 16380
rect 12348 16046 12350 16098
rect 12402 16046 12404 16098
rect 12348 16034 12404 16046
rect 12460 20018 12516 21196
rect 12572 21186 12628 21196
rect 12684 21140 12740 24444
rect 12796 23154 12852 24780
rect 13020 24742 13076 24780
rect 12908 24722 12964 24734
rect 12908 24670 12910 24722
rect 12962 24670 12964 24722
rect 12908 24276 12964 24670
rect 12908 23826 12964 24220
rect 13356 24276 13412 26908
rect 13468 26962 13524 26974
rect 13468 26910 13470 26962
rect 13522 26910 13524 26962
rect 13468 26516 13524 26910
rect 13468 26450 13524 26460
rect 13580 26962 13636 26974
rect 13580 26910 13582 26962
rect 13634 26910 13636 26962
rect 13580 26292 13636 26910
rect 13692 26964 13748 27002
rect 13692 26898 13748 26908
rect 13580 26226 13636 26236
rect 13804 26290 13860 27244
rect 13916 26740 13972 28140
rect 14028 27860 14084 27870
rect 14028 27634 14084 27804
rect 14028 27582 14030 27634
rect 14082 27582 14084 27634
rect 14028 27524 14084 27582
rect 14028 27458 14084 27468
rect 13916 26674 13972 26684
rect 14028 27186 14084 27198
rect 14028 27134 14030 27186
rect 14082 27134 14084 27186
rect 14028 27074 14084 27134
rect 14028 27022 14030 27074
rect 14082 27022 14084 27074
rect 13804 26238 13806 26290
rect 13858 26238 13860 26290
rect 13804 26226 13860 26238
rect 13916 26516 13972 26526
rect 13468 26180 13524 26190
rect 13468 26086 13524 26124
rect 13692 26066 13748 26078
rect 13916 26068 13972 26460
rect 13692 26014 13694 26066
rect 13746 26014 13748 26066
rect 13692 25956 13748 26014
rect 13692 25890 13748 25900
rect 13804 26012 13972 26068
rect 13804 25620 13860 26012
rect 13580 25282 13636 25294
rect 13580 25230 13582 25282
rect 13634 25230 13636 25282
rect 13580 25060 13636 25230
rect 13804 25060 13860 25564
rect 13916 25508 13972 25518
rect 13916 25414 13972 25452
rect 13580 24994 13636 25004
rect 13692 25004 13860 25060
rect 13468 24948 13524 24958
rect 13468 24722 13524 24892
rect 13468 24670 13470 24722
rect 13522 24670 13524 24722
rect 13468 24658 13524 24670
rect 13356 24210 13412 24220
rect 12908 23774 12910 23826
rect 12962 23774 12964 23826
rect 12908 23762 12964 23774
rect 12796 23102 12798 23154
rect 12850 23102 12852 23154
rect 12796 23090 12852 23102
rect 13468 22258 13524 22270
rect 13468 22206 13470 22258
rect 13522 22206 13524 22258
rect 13468 21924 13524 22206
rect 13468 21858 13524 21868
rect 13132 21588 13188 21598
rect 12684 21074 12740 21084
rect 12908 21474 12964 21486
rect 12908 21422 12910 21474
rect 12962 21422 12964 21474
rect 12908 20916 12964 21422
rect 12460 19966 12462 20018
rect 12514 19966 12516 20018
rect 12012 15374 12014 15426
rect 12066 15374 12068 15426
rect 12012 15362 12068 15374
rect 11788 15262 11790 15314
rect 11842 15262 11844 15314
rect 11788 15250 11844 15262
rect 11900 15202 11956 15214
rect 11900 15150 11902 15202
rect 11954 15150 11956 15202
rect 11788 15092 11844 15102
rect 11676 14532 11732 14542
rect 11788 14532 11844 15036
rect 11676 14530 11844 14532
rect 11676 14478 11678 14530
rect 11730 14478 11844 14530
rect 11676 14476 11844 14478
rect 11676 14466 11732 14476
rect 11452 14420 11508 14430
rect 11004 13356 11172 13412
rect 11228 14418 11508 14420
rect 11228 14366 11454 14418
rect 11506 14366 11508 14418
rect 11228 14364 11508 14366
rect 11228 13972 11284 14364
rect 11452 14354 11508 14364
rect 10780 12068 10836 12078
rect 10780 11974 10836 12012
rect 10668 11732 10948 11788
rect 10444 11666 10500 11676
rect 10108 11106 10164 11116
rect 10220 11396 10276 11406
rect 10220 10722 10276 11340
rect 10556 11394 10612 11406
rect 10556 11342 10558 11394
rect 10610 11342 10612 11394
rect 10556 10948 10612 11342
rect 10556 10882 10612 10892
rect 10220 10670 10222 10722
rect 10274 10670 10276 10722
rect 10220 10658 10276 10670
rect 10444 10836 10500 10846
rect 10444 10610 10500 10780
rect 10444 10558 10446 10610
rect 10498 10558 10500 10610
rect 10444 10546 10500 10558
rect 10556 10500 10612 10510
rect 10556 10406 10612 10444
rect 9772 9774 9774 9826
rect 9826 9774 9828 9826
rect 9772 9762 9828 9774
rect 10332 9828 10388 9838
rect 10332 9734 10388 9772
rect 10892 9826 10948 11732
rect 10892 9774 10894 9826
rect 10946 9774 10948 9826
rect 10892 9762 10948 9774
rect 9996 9604 10052 9614
rect 9884 9602 10052 9604
rect 9884 9550 9998 9602
rect 10050 9550 10052 9602
rect 9884 9548 10052 9550
rect 9884 8260 9940 9548
rect 9996 9538 10052 9548
rect 9996 9380 10052 9390
rect 11004 9380 11060 13356
rect 11228 13300 11284 13916
rect 11788 13972 11844 13982
rect 11340 13748 11396 13758
rect 11340 13654 11396 13692
rect 11116 13244 11284 13300
rect 11116 12178 11172 13244
rect 11340 12962 11396 12974
rect 11340 12910 11342 12962
rect 11394 12910 11396 12962
rect 11228 12850 11284 12862
rect 11228 12798 11230 12850
rect 11282 12798 11284 12850
rect 11228 12404 11284 12798
rect 11228 12338 11284 12348
rect 11116 12126 11118 12178
rect 11170 12126 11172 12178
rect 11116 12114 11172 12126
rect 11340 12292 11396 12910
rect 11564 12292 11620 12302
rect 11340 12290 11620 12292
rect 11340 12238 11566 12290
rect 11618 12238 11620 12290
rect 11340 12236 11620 12238
rect 11340 12180 11396 12236
rect 11340 12114 11396 12124
rect 11228 11620 11284 11630
rect 11228 11170 11284 11564
rect 11228 11118 11230 11170
rect 11282 11118 11284 11170
rect 11116 9380 11172 9390
rect 11004 9324 11116 9380
rect 9996 9266 10052 9324
rect 11116 9314 11172 9324
rect 9996 9214 9998 9266
rect 10050 9214 10052 9266
rect 9996 9202 10052 9214
rect 10892 9268 10948 9278
rect 10444 9044 10500 9054
rect 10444 8950 10500 8988
rect 10892 8370 10948 9212
rect 10892 8318 10894 8370
rect 10946 8318 10948 8370
rect 10892 8306 10948 8318
rect 9884 8194 9940 8204
rect 9884 7700 9940 7710
rect 9660 7698 10276 7700
rect 9660 7646 9886 7698
rect 9938 7646 10276 7698
rect 9660 7644 10276 7646
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 9884 6804 9940 7644
rect 10220 7474 10276 7644
rect 10220 7422 10222 7474
rect 10274 7422 10276 7474
rect 10220 7410 10276 7422
rect 10668 7474 10724 7486
rect 10668 7422 10670 7474
rect 10722 7422 10724 7474
rect 10668 7028 10724 7422
rect 11004 7476 11060 7486
rect 11004 7382 11060 7420
rect 10892 7028 10948 7038
rect 10668 6972 10892 7028
rect 10892 6962 10948 6972
rect 9884 6710 9940 6748
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 11228 3388 11284 11118
rect 11452 10612 11508 10622
rect 11452 10518 11508 10556
rect 11564 9714 11620 12236
rect 11788 12290 11844 13916
rect 11900 13748 11956 15150
rect 12124 14642 12180 14654
rect 12124 14590 12126 14642
rect 12178 14590 12180 14642
rect 11900 13682 11956 13692
rect 12012 14418 12068 14430
rect 12012 14366 12014 14418
rect 12066 14366 12068 14418
rect 11788 12238 11790 12290
rect 11842 12238 11844 12290
rect 11788 12226 11844 12238
rect 11900 12962 11956 12974
rect 11900 12910 11902 12962
rect 11954 12910 11956 12962
rect 11900 12292 11956 12910
rect 12012 12516 12068 14366
rect 12124 14420 12180 14590
rect 12124 14354 12180 14364
rect 12012 12450 12068 12460
rect 12124 13074 12180 13086
rect 12124 13022 12126 13074
rect 12178 13022 12180 13074
rect 12124 12292 12180 13022
rect 12460 13076 12516 19966
rect 12572 20860 12964 20916
rect 12572 19796 12628 20860
rect 12684 20690 12740 20702
rect 12684 20638 12686 20690
rect 12738 20638 12740 20690
rect 12684 20244 12740 20638
rect 12684 20178 12740 20188
rect 12796 20578 12852 20590
rect 13020 20580 13076 20590
rect 12796 20526 12798 20578
rect 12850 20526 12852 20578
rect 12796 19908 12852 20526
rect 12908 20578 13076 20580
rect 12908 20526 13022 20578
rect 13074 20526 13076 20578
rect 12908 20524 13076 20526
rect 12908 20020 12964 20524
rect 13020 20514 13076 20524
rect 12908 19954 12964 19964
rect 13020 20018 13076 20030
rect 13020 19966 13022 20018
rect 13074 19966 13076 20018
rect 12796 19842 12852 19852
rect 12572 19012 12628 19740
rect 12572 18946 12628 18956
rect 13020 18900 13076 19966
rect 13020 18834 13076 18844
rect 13132 18452 13188 21532
rect 13692 21588 13748 25004
rect 13916 24164 13972 24174
rect 13916 23716 13972 24108
rect 13916 23622 13972 23660
rect 13916 23380 13972 23390
rect 13916 22930 13972 23324
rect 13916 22878 13918 22930
rect 13970 22878 13972 22930
rect 13692 21522 13748 21532
rect 13804 22596 13860 22606
rect 13132 18386 13188 18396
rect 13356 21476 13412 21486
rect 13356 18900 13412 21420
rect 13692 20802 13748 20814
rect 13692 20750 13694 20802
rect 13746 20750 13748 20802
rect 13468 20692 13524 20702
rect 13468 20598 13524 20636
rect 13692 20580 13748 20750
rect 13692 20514 13748 20524
rect 13804 20244 13860 22540
rect 13916 22260 13972 22878
rect 13916 22194 13972 22204
rect 13580 20188 13860 20244
rect 13916 20914 13972 20926
rect 13916 20862 13918 20914
rect 13970 20862 13972 20914
rect 13356 18450 13412 18844
rect 13468 20018 13524 20030
rect 13468 19966 13470 20018
rect 13522 19966 13524 20018
rect 13468 19572 13524 19966
rect 13468 18676 13524 19516
rect 13580 19346 13636 20188
rect 13692 20020 13748 20030
rect 13692 19926 13748 19964
rect 13580 19294 13582 19346
rect 13634 19294 13636 19346
rect 13580 19282 13636 19294
rect 13916 19796 13972 20862
rect 13468 18610 13524 18620
rect 13356 18398 13358 18450
rect 13410 18398 13412 18450
rect 13356 18386 13412 18398
rect 13692 18452 13748 18462
rect 13692 18358 13748 18396
rect 13580 18340 13636 18350
rect 13580 17666 13636 18284
rect 13580 17614 13582 17666
rect 13634 17614 13636 17666
rect 12908 17556 12964 17566
rect 12908 17462 12964 17500
rect 13580 16884 13636 17614
rect 13916 17554 13972 19740
rect 14028 19124 14084 27022
rect 14140 25844 14196 29708
rect 14364 29428 14420 29438
rect 14364 29334 14420 29372
rect 15372 29428 15428 29438
rect 14924 29314 14980 29326
rect 14924 29262 14926 29314
rect 14978 29262 14980 29314
rect 14700 28644 14756 28654
rect 14700 28550 14756 28588
rect 14252 28418 14308 28430
rect 14252 28366 14254 28418
rect 14306 28366 14308 28418
rect 14252 27298 14308 28366
rect 14364 27748 14420 27758
rect 14364 27654 14420 27692
rect 14924 27412 14980 29262
rect 15372 28868 15428 29372
rect 15596 29428 15652 29438
rect 15596 29334 15652 29372
rect 16044 29314 16100 29326
rect 16044 29262 16046 29314
rect 16098 29262 16100 29314
rect 15372 28812 15652 28868
rect 15036 28754 15092 28766
rect 15036 28702 15038 28754
rect 15090 28702 15092 28754
rect 15036 27972 15092 28702
rect 15484 28644 15540 28654
rect 15484 28550 15540 28588
rect 15596 28532 15652 28812
rect 16044 28756 16100 29262
rect 16716 29316 16772 29326
rect 16716 29222 16772 29260
rect 16044 28690 16100 28700
rect 16380 28756 16436 28766
rect 16380 28642 16436 28700
rect 16380 28590 16382 28642
rect 16434 28590 16436 28642
rect 16380 28578 16436 28590
rect 16044 28532 16100 28542
rect 15596 28082 15652 28476
rect 15596 28030 15598 28082
rect 15650 28030 15652 28082
rect 15596 28018 15652 28030
rect 15932 28530 16100 28532
rect 15932 28478 16046 28530
rect 16098 28478 16100 28530
rect 15932 28476 16100 28478
rect 15148 27972 15204 27982
rect 15036 27916 15148 27972
rect 15148 27906 15204 27916
rect 14252 27246 14254 27298
rect 14306 27246 14308 27298
rect 14252 27188 14308 27246
rect 14252 27122 14308 27132
rect 14588 27356 14980 27412
rect 15148 27746 15204 27758
rect 15148 27694 15150 27746
rect 15202 27694 15204 27746
rect 14476 27074 14532 27086
rect 14476 27022 14478 27074
rect 14530 27022 14532 27074
rect 14252 26740 14308 26750
rect 14252 26290 14308 26684
rect 14252 26238 14254 26290
rect 14306 26238 14308 26290
rect 14252 26068 14308 26238
rect 14252 26002 14308 26012
rect 14140 25732 14196 25788
rect 14476 25732 14532 27022
rect 14588 26908 14644 27356
rect 14700 27188 14756 27198
rect 14700 27076 14756 27132
rect 14924 27076 14980 27086
rect 14700 27074 14980 27076
rect 14700 27022 14926 27074
rect 14978 27022 14980 27074
rect 14700 27020 14980 27022
rect 14924 27010 14980 27020
rect 14588 26852 15092 26908
rect 15036 26516 15092 26852
rect 14140 25676 14420 25732
rect 14364 25620 14420 25676
rect 14364 25554 14420 25564
rect 14140 25506 14196 25518
rect 14140 25454 14142 25506
rect 14194 25454 14196 25506
rect 14140 24948 14196 25454
rect 14140 24882 14196 24892
rect 14252 25508 14308 25518
rect 14252 23380 14308 25452
rect 14252 23314 14308 23324
rect 14364 24612 14420 24622
rect 14364 23940 14420 24556
rect 14476 24164 14532 25676
rect 14588 26460 15092 26516
rect 14588 25060 14644 26460
rect 14700 26292 14756 26302
rect 15148 26292 15204 27694
rect 15708 27076 15764 27114
rect 15708 27010 15764 27020
rect 15932 26908 15988 28476
rect 16044 28466 16100 28476
rect 16716 28532 16772 28542
rect 16716 28438 16772 28476
rect 16268 27972 16324 27982
rect 16324 27916 16436 27972
rect 16268 27878 16324 27916
rect 16268 27300 16324 27310
rect 15708 26852 15988 26908
rect 16044 26962 16100 26974
rect 16044 26910 16046 26962
rect 16098 26910 16100 26962
rect 15372 26628 15428 26638
rect 14700 26290 15204 26292
rect 14700 26238 14702 26290
rect 14754 26238 15204 26290
rect 14700 26236 15204 26238
rect 15260 26292 15316 26302
rect 14700 26226 14756 26236
rect 14812 25956 14868 25966
rect 14812 25620 14868 25900
rect 14812 25554 14868 25564
rect 14812 25172 14868 25182
rect 14700 25060 14756 25070
rect 14588 25004 14700 25060
rect 14700 24994 14756 25004
rect 14476 24108 14644 24164
rect 14476 23940 14532 23950
rect 14364 23938 14532 23940
rect 14364 23886 14478 23938
rect 14530 23886 14532 23938
rect 14364 23884 14532 23886
rect 14140 23154 14196 23166
rect 14140 23102 14142 23154
rect 14194 23102 14196 23154
rect 14140 22370 14196 23102
rect 14140 22318 14142 22370
rect 14194 22318 14196 22370
rect 14140 21700 14196 22318
rect 14252 21700 14308 21710
rect 14196 21698 14308 21700
rect 14196 21646 14254 21698
rect 14306 21646 14308 21698
rect 14196 21644 14308 21646
rect 14140 21606 14196 21644
rect 14252 21634 14308 21644
rect 14140 20692 14196 20702
rect 14140 19346 14196 20636
rect 14140 19294 14142 19346
rect 14194 19294 14196 19346
rect 14140 19282 14196 19294
rect 14252 19236 14308 19246
rect 14252 19142 14308 19180
rect 14028 19058 14084 19068
rect 14364 19012 14420 23884
rect 14476 23874 14532 23884
rect 14588 23828 14644 24108
rect 14812 23938 14868 25116
rect 15036 25172 15092 26236
rect 15260 26198 15316 26236
rect 15372 25956 15428 26572
rect 15596 26402 15652 26414
rect 15596 26350 15598 26402
rect 15650 26350 15652 26402
rect 15596 26068 15652 26350
rect 15596 26002 15652 26012
rect 15372 25844 15428 25900
rect 15260 25788 15428 25844
rect 15260 25506 15316 25788
rect 15260 25454 15262 25506
rect 15314 25454 15316 25506
rect 15260 25442 15316 25454
rect 15372 25618 15428 25630
rect 15372 25566 15374 25618
rect 15426 25566 15428 25618
rect 15372 25508 15428 25566
rect 15372 25442 15428 25452
rect 15036 25106 15092 25116
rect 15484 25396 15540 25406
rect 15708 25396 15764 26852
rect 16044 25620 16100 26910
rect 16268 26964 16324 27244
rect 16268 26898 16324 26908
rect 16268 26514 16324 26526
rect 16268 26462 16270 26514
rect 16322 26462 16324 26514
rect 16156 26292 16212 26302
rect 16156 26198 16212 26236
rect 16268 25844 16324 26462
rect 16268 25778 16324 25788
rect 16044 25564 16212 25620
rect 15932 25508 15988 25518
rect 15932 25414 15988 25452
rect 15484 25394 15764 25396
rect 15484 25342 15486 25394
rect 15538 25342 15764 25394
rect 15484 25340 15764 25342
rect 14924 24834 14980 24846
rect 14924 24782 14926 24834
rect 14978 24782 14980 24834
rect 14924 24276 14980 24782
rect 15484 24612 15540 25340
rect 15820 25172 15876 25182
rect 14924 24210 14980 24220
rect 15148 24556 15540 24612
rect 15708 25060 15764 25070
rect 14812 23886 14814 23938
rect 14866 23886 14868 23938
rect 14700 23828 14756 23838
rect 14588 23772 14700 23828
rect 14588 20916 14644 20926
rect 14476 20020 14532 20030
rect 14476 19348 14532 19964
rect 14476 19282 14532 19292
rect 13916 17502 13918 17554
rect 13970 17502 13972 17554
rect 13916 17490 13972 17502
rect 14140 18956 14420 19012
rect 14140 17332 14196 18956
rect 14588 18450 14644 20860
rect 14588 18398 14590 18450
rect 14642 18398 14644 18450
rect 13580 16818 13636 16828
rect 13804 17276 14196 17332
rect 14252 18338 14308 18350
rect 14588 18340 14644 18398
rect 14252 18286 14254 18338
rect 14306 18286 14308 18338
rect 13468 16772 13524 16782
rect 13356 16716 13468 16772
rect 13356 16212 13412 16716
rect 13468 16678 13524 16716
rect 13356 16146 13412 16156
rect 13692 16548 13748 16558
rect 13580 16100 13636 16110
rect 12572 15764 12628 15774
rect 12572 15314 12628 15708
rect 13580 15764 13636 16044
rect 13580 15698 13636 15708
rect 13692 15986 13748 16492
rect 13692 15934 13694 15986
rect 13746 15934 13748 15986
rect 12572 15262 12574 15314
rect 12626 15262 12628 15314
rect 12572 15250 12628 15262
rect 13132 15540 13188 15550
rect 12908 14980 12964 14990
rect 12572 14532 12628 14542
rect 12572 14438 12628 14476
rect 12684 14420 12740 14430
rect 12684 13746 12740 14364
rect 12684 13694 12686 13746
rect 12738 13694 12740 13746
rect 12684 13682 12740 13694
rect 12908 13076 12964 14924
rect 13132 13746 13188 15484
rect 13692 15316 13748 15934
rect 13692 15250 13748 15260
rect 13356 15202 13412 15214
rect 13356 15150 13358 15202
rect 13410 15150 13412 15202
rect 13356 15148 13412 15150
rect 13356 15092 13636 15148
rect 13132 13694 13134 13746
rect 13186 13694 13188 13746
rect 13132 13682 13188 13694
rect 13468 14644 13524 14654
rect 13244 13524 13300 13534
rect 12460 13020 12628 13076
rect 11900 12226 11956 12236
rect 12012 12236 12180 12292
rect 12348 12852 12404 12862
rect 11676 12180 11732 12190
rect 11676 12068 11732 12124
rect 11676 12012 11844 12068
rect 11564 9662 11566 9714
rect 11618 9662 11620 9714
rect 11340 8932 11396 8942
rect 11340 8838 11396 8876
rect 11340 8708 11396 8718
rect 11340 8370 11396 8652
rect 11340 8318 11342 8370
rect 11394 8318 11396 8370
rect 11340 8306 11396 8318
rect 11564 8258 11620 9662
rect 11676 10052 11732 10062
rect 11676 9826 11732 9996
rect 11676 9774 11678 9826
rect 11730 9774 11732 9826
rect 11676 8932 11732 9774
rect 11788 9266 11844 12012
rect 11900 12066 11956 12078
rect 11900 12014 11902 12066
rect 11954 12014 11956 12066
rect 11900 11620 11956 12014
rect 11900 11554 11956 11564
rect 11900 11396 11956 11406
rect 12012 11396 12068 12236
rect 12348 12178 12404 12796
rect 12348 12126 12350 12178
rect 12402 12126 12404 12178
rect 12348 12114 12404 12126
rect 12460 12850 12516 12862
rect 12460 12798 12462 12850
rect 12514 12798 12516 12850
rect 11956 11340 12068 11396
rect 11900 11302 11956 11340
rect 12348 11284 12404 11294
rect 12236 11228 12348 11284
rect 12236 10388 12292 11228
rect 12348 11190 12404 11228
rect 12348 10612 12404 10622
rect 12460 10612 12516 12798
rect 12404 10556 12516 10612
rect 12572 10836 12628 13020
rect 12908 12982 12964 13020
rect 13132 13522 13300 13524
rect 13132 13470 13246 13522
rect 13298 13470 13300 13522
rect 13132 13468 13300 13470
rect 12796 11732 12852 11742
rect 12796 11394 12852 11676
rect 12796 11342 12798 11394
rect 12850 11342 12852 11394
rect 12796 11330 12852 11342
rect 12908 11172 12964 11182
rect 12348 10546 12404 10556
rect 12236 10332 12404 10388
rect 12236 9828 12292 9838
rect 12124 9604 12180 9614
rect 11788 9214 11790 9266
rect 11842 9214 11844 9266
rect 11788 9202 11844 9214
rect 11900 9602 12180 9604
rect 11900 9550 12126 9602
rect 12178 9550 12180 9602
rect 11900 9548 12180 9550
rect 11676 8866 11732 8876
rect 11900 8260 11956 9548
rect 12124 9538 12180 9548
rect 11564 8206 11566 8258
rect 11618 8206 11620 8258
rect 11564 8194 11620 8206
rect 11788 8204 11956 8260
rect 12124 9156 12180 9166
rect 12236 9156 12292 9772
rect 12124 9154 12292 9156
rect 12124 9102 12126 9154
rect 12178 9102 12292 9154
rect 12124 9100 12292 9102
rect 11676 7476 11732 7486
rect 11676 6690 11732 7420
rect 11676 6638 11678 6690
rect 11730 6638 11732 6690
rect 11676 6626 11732 6638
rect 11340 6580 11396 6590
rect 11340 6486 11396 6524
rect 4732 3332 4788 3342
rect 4732 800 4788 3276
rect 5516 3332 5572 3342
rect 9660 3332 9716 3342
rect 11228 3332 11620 3388
rect 5516 3238 5572 3276
rect 9436 3330 9716 3332
rect 9436 3278 9662 3330
rect 9714 3278 9716 3330
rect 9436 3276 9716 3278
rect 9436 800 9492 3276
rect 9660 3266 9716 3276
rect 11564 3266 11620 3276
rect 11788 2884 11844 8204
rect 12012 8148 12068 8158
rect 11900 8034 11956 8046
rect 11900 7982 11902 8034
rect 11954 7982 11956 8034
rect 11900 6692 11956 7982
rect 12012 7474 12068 8092
rect 12012 7422 12014 7474
rect 12066 7422 12068 7474
rect 12012 7410 12068 7422
rect 12124 7028 12180 9100
rect 12236 8932 12292 8942
rect 12236 8034 12292 8876
rect 12348 8708 12404 10332
rect 12572 9042 12628 10780
rect 12796 10948 12852 10958
rect 12796 10610 12852 10892
rect 12908 10836 12964 11116
rect 12908 10770 12964 10780
rect 12796 10558 12798 10610
rect 12850 10558 12852 10610
rect 12796 9940 12852 10558
rect 12796 9874 12852 9884
rect 12572 8990 12574 9042
rect 12626 8990 12628 9042
rect 12572 8978 12628 8990
rect 13020 9602 13076 9614
rect 13020 9550 13022 9602
rect 13074 9550 13076 9602
rect 12684 8932 12740 8942
rect 12684 8838 12740 8876
rect 12348 8642 12404 8652
rect 13020 8596 13076 9550
rect 13020 8530 13076 8540
rect 13132 8484 13188 13468
rect 13244 13458 13300 13468
rect 13244 13076 13300 13086
rect 13244 12402 13300 13020
rect 13244 12350 13246 12402
rect 13298 12350 13300 12402
rect 13244 12338 13300 12350
rect 13468 12178 13524 14588
rect 13580 14642 13636 15092
rect 13580 14590 13582 14642
rect 13634 14590 13636 14642
rect 13580 14578 13636 14590
rect 13692 14868 13748 14878
rect 13692 14530 13748 14812
rect 13692 14478 13694 14530
rect 13746 14478 13748 14530
rect 13692 14084 13748 14478
rect 13468 12126 13470 12178
rect 13522 12126 13524 12178
rect 13468 12114 13524 12126
rect 13580 14028 13692 14084
rect 13580 11508 13636 14028
rect 13692 14018 13748 14028
rect 13692 12740 13748 12750
rect 13692 12646 13748 12684
rect 13580 11452 13748 11508
rect 13692 11172 13748 11452
rect 13804 11396 13860 17276
rect 13916 16884 13972 16894
rect 13916 14418 13972 16828
rect 14028 15876 14084 15886
rect 14028 15782 14084 15820
rect 14140 15652 14196 15662
rect 14140 15314 14196 15596
rect 14252 15540 14308 18286
rect 14364 18284 14644 18340
rect 14700 18340 14756 23772
rect 14812 21586 14868 23886
rect 15148 23828 15204 24556
rect 15708 24276 15764 25004
rect 15820 24948 15876 25116
rect 16156 24948 16212 25564
rect 15820 24946 16212 24948
rect 15820 24894 16158 24946
rect 16210 24894 16212 24946
rect 15820 24892 16212 24894
rect 15820 24722 15876 24892
rect 16156 24882 16212 24892
rect 16268 25394 16324 25406
rect 16268 25342 16270 25394
rect 16322 25342 16324 25394
rect 16268 24948 16324 25342
rect 15820 24670 15822 24722
rect 15874 24670 15876 24722
rect 15820 24658 15876 24670
rect 15932 24276 15988 24286
rect 15708 24220 15932 24276
rect 15372 23938 15428 23950
rect 15372 23886 15374 23938
rect 15426 23886 15428 23938
rect 15148 23772 15316 23828
rect 14812 21534 14814 21586
rect 14866 21534 14868 21586
rect 14812 20132 14868 21534
rect 14812 20066 14868 20076
rect 14924 23154 14980 23166
rect 14924 23102 14926 23154
rect 14978 23102 14980 23154
rect 14924 21476 14980 23102
rect 15036 21476 15092 21486
rect 14924 21474 15092 21476
rect 14924 21422 15038 21474
rect 15090 21422 15092 21474
rect 14924 21420 15092 21422
rect 14812 19236 14868 19246
rect 14924 19236 14980 21420
rect 15036 21410 15092 21420
rect 15260 21252 15316 23772
rect 15372 21364 15428 23886
rect 15708 23940 15764 23950
rect 15708 23826 15764 23884
rect 15932 23938 15988 24220
rect 15932 23886 15934 23938
rect 15986 23886 15988 23938
rect 15932 23874 15988 23886
rect 16044 24052 16100 24062
rect 15708 23774 15710 23826
rect 15762 23774 15764 23826
rect 15708 23762 15764 23774
rect 15708 23042 15764 23054
rect 15708 22990 15710 23042
rect 15762 22990 15764 23042
rect 15372 21298 15428 21308
rect 15484 22930 15540 22942
rect 15484 22878 15486 22930
rect 15538 22878 15540 22930
rect 15036 21196 15316 21252
rect 15036 20916 15092 21196
rect 15036 20850 15092 20860
rect 15148 21028 15204 21038
rect 15484 21028 15540 22878
rect 15708 22708 15764 22990
rect 16044 22708 16100 23996
rect 16268 23492 16324 24892
rect 16268 23426 16324 23436
rect 16156 23044 16212 23054
rect 16156 22950 16212 22988
rect 16380 22930 16436 27916
rect 16828 27746 16884 27758
rect 16828 27694 16830 27746
rect 16882 27694 16884 27746
rect 16828 27412 16884 27694
rect 16828 27346 16884 27356
rect 16604 27188 16660 27198
rect 16604 27094 16660 27132
rect 16716 26292 16772 26302
rect 16492 25618 16548 25630
rect 16492 25566 16494 25618
rect 16546 25566 16548 25618
rect 16492 25284 16548 25566
rect 16492 25218 16548 25228
rect 16604 24612 16660 24622
rect 16604 24518 16660 24556
rect 16716 24388 16772 26236
rect 16828 26180 16884 26190
rect 16828 26086 16884 26124
rect 16604 24332 16772 24388
rect 17052 25506 17108 30492
rect 17500 29540 17556 30940
rect 17612 30212 17668 30222
rect 17836 30212 17892 30222
rect 17612 30210 17780 30212
rect 17612 30158 17614 30210
rect 17666 30158 17780 30210
rect 17612 30156 17780 30158
rect 17612 30146 17668 30156
rect 17500 29474 17556 29484
rect 17724 29652 17780 30156
rect 17836 30210 18116 30212
rect 17836 30158 17838 30210
rect 17890 30158 18116 30210
rect 17836 30156 18116 30158
rect 17836 30146 17892 30156
rect 17612 29428 17668 29438
rect 17612 28644 17668 29372
rect 17724 29204 17780 29596
rect 18060 29988 18116 30156
rect 18396 30098 18452 31500
rect 18956 31554 19124 31556
rect 18956 31502 18958 31554
rect 19010 31502 19124 31554
rect 18956 31500 19124 31502
rect 19180 32900 19236 32910
rect 18956 31220 19012 31500
rect 18956 31154 19012 31164
rect 19180 31220 19236 32844
rect 19180 31154 19236 31164
rect 19292 31668 19348 31678
rect 19404 31668 19460 34076
rect 19516 34038 19572 34076
rect 19740 34130 19796 34142
rect 19740 34078 19742 34130
rect 19794 34078 19796 34130
rect 19516 33796 19572 33806
rect 19740 33796 19796 34078
rect 19852 34130 19908 34300
rect 20524 34244 20580 36876
rect 20636 34804 20692 37212
rect 20748 37202 20804 37212
rect 20972 37268 21028 43486
rect 21420 43316 21476 46396
rect 21532 46386 21588 46396
rect 21644 45780 21700 45790
rect 21532 45666 21588 45678
rect 21532 45614 21534 45666
rect 21586 45614 21588 45666
rect 21532 45444 21588 45614
rect 21532 45378 21588 45388
rect 21644 44772 21700 45724
rect 21756 45330 21812 48188
rect 21868 48132 21924 51548
rect 21980 50428 22036 54236
rect 22092 54226 22148 54236
rect 22428 53620 22484 53630
rect 22428 53526 22484 53564
rect 22540 53060 22596 54460
rect 22764 53170 22820 55580
rect 22764 53118 22766 53170
rect 22818 53118 22820 53170
rect 22764 53106 22820 53118
rect 22540 52966 22596 53004
rect 22540 52164 22596 52174
rect 22540 52070 22596 52108
rect 22876 52052 22932 57372
rect 22988 57362 23044 57372
rect 24780 56420 24836 56430
rect 23324 56308 23380 56318
rect 23324 56214 23380 56252
rect 24668 56196 24724 56206
rect 24668 56102 24724 56140
rect 23548 56084 23604 56094
rect 23100 55972 23156 55982
rect 23100 55970 23268 55972
rect 23100 55918 23102 55970
rect 23154 55918 23268 55970
rect 23100 55916 23268 55918
rect 23100 55906 23156 55916
rect 23212 55524 23268 55916
rect 23100 55074 23156 55086
rect 23100 55022 23102 55074
rect 23154 55022 23156 55074
rect 23100 53844 23156 55022
rect 23100 53778 23156 53788
rect 22764 51996 22932 52052
rect 22988 53620 23044 53630
rect 22988 52276 23044 53564
rect 23212 53058 23268 55468
rect 23548 55188 23604 56028
rect 24556 56082 24612 56094
rect 24556 56030 24558 56082
rect 24610 56030 24612 56082
rect 24556 55860 24612 56030
rect 24556 55794 24612 55804
rect 24668 55858 24724 55870
rect 24668 55806 24670 55858
rect 24722 55806 24724 55858
rect 24332 55412 24388 55422
rect 24332 55318 24388 55356
rect 23548 54404 23604 55132
rect 23772 55298 23828 55310
rect 23996 55300 24052 55310
rect 23772 55246 23774 55298
rect 23826 55246 23828 55298
rect 23772 54852 23828 55246
rect 23772 54786 23828 54796
rect 23884 55298 24052 55300
rect 23884 55246 23998 55298
rect 24050 55246 24052 55298
rect 23884 55244 24052 55246
rect 23548 54338 23604 54348
rect 23660 54628 23716 54638
rect 23884 54628 23940 55244
rect 23996 55234 24052 55244
rect 23660 54626 23940 54628
rect 23660 54574 23662 54626
rect 23714 54574 23940 54626
rect 23660 54572 23940 54574
rect 23996 54626 24052 54638
rect 23996 54574 23998 54626
rect 24050 54574 24052 54626
rect 23436 53844 23492 53854
rect 23492 53788 23604 53844
rect 23436 53778 23492 53788
rect 23212 53006 23214 53058
rect 23266 53006 23268 53058
rect 23212 52994 23268 53006
rect 23436 53618 23492 53630
rect 23436 53566 23438 53618
rect 23490 53566 23492 53618
rect 22316 51938 22372 51950
rect 22316 51886 22318 51938
rect 22370 51886 22372 51938
rect 22316 51492 22372 51886
rect 22316 51426 22372 51436
rect 22540 51380 22596 51390
rect 22428 51378 22596 51380
rect 22428 51326 22542 51378
rect 22594 51326 22596 51378
rect 22428 51324 22596 51326
rect 22204 51154 22260 51166
rect 22204 51102 22206 51154
rect 22258 51102 22260 51154
rect 22204 50596 22260 51102
rect 22204 50530 22260 50540
rect 22428 50428 22484 51324
rect 22540 51314 22596 51324
rect 22540 51156 22596 51166
rect 22540 51062 22596 51100
rect 21980 50372 22148 50428
rect 22428 50372 22596 50428
rect 22092 49700 22148 50372
rect 22148 49644 22372 49700
rect 22092 49634 22148 49644
rect 22316 49026 22372 49644
rect 22316 48974 22318 49026
rect 22370 48974 22372 49026
rect 22316 48962 22372 48974
rect 22428 49138 22484 49150
rect 22428 49086 22430 49138
rect 22482 49086 22484 49138
rect 21868 48066 21924 48076
rect 22316 48242 22372 48254
rect 22316 48190 22318 48242
rect 22370 48190 22372 48242
rect 22316 47684 22372 48190
rect 22316 47618 22372 47628
rect 22428 47570 22484 49086
rect 22428 47518 22430 47570
rect 22482 47518 22484 47570
rect 22428 47506 22484 47518
rect 22316 47346 22372 47358
rect 22316 47294 22318 47346
rect 22370 47294 22372 47346
rect 21868 47234 21924 47246
rect 21868 47182 21870 47234
rect 21922 47182 21924 47234
rect 21868 47012 21924 47182
rect 21868 46946 21924 46956
rect 22204 46676 22260 46686
rect 21868 46674 22260 46676
rect 21868 46622 22206 46674
rect 22258 46622 22260 46674
rect 21868 46620 22260 46622
rect 21868 46562 21924 46620
rect 22204 46610 22260 46620
rect 21868 46510 21870 46562
rect 21922 46510 21924 46562
rect 21868 46498 21924 46510
rect 21868 46228 21924 46238
rect 21868 45890 21924 46172
rect 21868 45838 21870 45890
rect 21922 45838 21924 45890
rect 21868 45826 21924 45838
rect 22092 46116 22148 46126
rect 21756 45278 21758 45330
rect 21810 45278 21812 45330
rect 21756 45266 21812 45278
rect 21980 45778 22036 45790
rect 21980 45726 21982 45778
rect 22034 45726 22036 45778
rect 21644 44716 21812 44772
rect 21644 43428 21700 43438
rect 21644 43334 21700 43372
rect 21420 43250 21476 43260
rect 21756 43316 21812 44716
rect 21868 44324 21924 44334
rect 21868 44230 21924 44268
rect 21756 43250 21812 43260
rect 21868 44100 21924 44110
rect 21868 43538 21924 44044
rect 21868 43486 21870 43538
rect 21922 43486 21924 43538
rect 21868 42980 21924 43486
rect 21980 43204 22036 45726
rect 21980 43138 22036 43148
rect 22092 44994 22148 46060
rect 22204 45556 22260 45566
rect 22316 45556 22372 47294
rect 22540 47124 22596 50372
rect 22764 50036 22820 51996
rect 22988 51604 23044 52220
rect 23324 52836 23380 52846
rect 23436 52836 23492 53566
rect 23548 53396 23604 53788
rect 23548 53058 23604 53340
rect 23548 53006 23550 53058
rect 23602 53006 23604 53058
rect 23548 52994 23604 53006
rect 23436 52780 23604 52836
rect 23324 52274 23380 52780
rect 23324 52222 23326 52274
rect 23378 52222 23380 52274
rect 22988 51602 23156 51604
rect 22988 51550 22990 51602
rect 23042 51550 23156 51602
rect 22988 51548 23156 51550
rect 22988 51538 23044 51548
rect 22876 51380 22932 51390
rect 22876 51286 22932 51324
rect 22988 51154 23044 51166
rect 22988 51102 22990 51154
rect 23042 51102 23044 51154
rect 22988 50372 23044 51102
rect 22988 50306 23044 50316
rect 22876 50036 22932 50046
rect 22764 50034 22932 50036
rect 22764 49982 22878 50034
rect 22930 49982 22932 50034
rect 22764 49980 22932 49982
rect 22876 49970 22932 49980
rect 22988 50036 23044 50046
rect 22764 49812 22820 49822
rect 22764 49718 22820 49756
rect 22988 48914 23044 49980
rect 23100 49924 23156 51548
rect 23100 49858 23156 49868
rect 23324 49476 23380 52222
rect 23548 51380 23604 52780
rect 23660 52612 23716 54572
rect 23884 54404 23940 54414
rect 23884 53844 23940 54348
rect 23660 52546 23716 52556
rect 23772 53788 23940 53844
rect 23772 52274 23828 53788
rect 23772 52222 23774 52274
rect 23826 52222 23828 52274
rect 23548 51314 23604 51324
rect 23660 52164 23716 52174
rect 23324 49410 23380 49420
rect 23548 51156 23604 51166
rect 22988 48862 22990 48914
rect 23042 48862 23044 48914
rect 22988 48850 23044 48862
rect 23324 49028 23380 49038
rect 22764 48804 22820 48814
rect 22764 47460 22820 48748
rect 22764 47366 22820 47404
rect 22876 48692 22932 48702
rect 22876 48242 22932 48636
rect 23324 48466 23380 48972
rect 23548 49026 23604 51100
rect 23660 50594 23716 52108
rect 23772 50708 23828 52222
rect 23996 52164 24052 54574
rect 24556 54516 24612 54526
rect 24556 54422 24612 54460
rect 24668 54404 24724 55806
rect 24780 55860 24836 56364
rect 24780 55794 24836 55804
rect 24220 54292 24276 54302
rect 24220 54198 24276 54236
rect 24108 53732 24164 53742
rect 24108 53638 24164 53676
rect 24332 53508 24388 53518
rect 24668 53508 24724 54348
rect 24220 53506 24388 53508
rect 24220 53454 24334 53506
rect 24386 53454 24388 53506
rect 24220 53452 24388 53454
rect 23996 52098 24052 52108
rect 24108 52834 24164 52846
rect 24108 52782 24110 52834
rect 24162 52782 24164 52834
rect 24108 51716 24164 52782
rect 24220 52162 24276 53452
rect 24332 53442 24388 53452
rect 24556 53452 24668 53508
rect 24332 53172 24388 53182
rect 24332 53078 24388 53116
rect 24220 52110 24222 52162
rect 24274 52110 24276 52162
rect 24220 52098 24276 52110
rect 24444 53060 24500 53070
rect 24444 52162 24500 53004
rect 24444 52110 24446 52162
rect 24498 52110 24500 52162
rect 24444 52098 24500 52110
rect 24556 51940 24612 53452
rect 24668 53442 24724 53452
rect 24892 54852 24948 54862
rect 24668 53060 24724 53070
rect 24668 52966 24724 53004
rect 23996 51660 24108 51716
rect 23884 51266 23940 51278
rect 23884 51214 23886 51266
rect 23938 51214 23940 51266
rect 23884 50820 23940 51214
rect 23884 50754 23940 50764
rect 23772 50642 23828 50652
rect 23660 50542 23662 50594
rect 23714 50542 23716 50594
rect 23660 50530 23716 50542
rect 23996 50596 24052 51660
rect 24108 51650 24164 51660
rect 24220 51884 24612 51940
rect 24780 52612 24836 52622
rect 24220 51380 24276 51884
rect 24220 51286 24276 51324
rect 23996 50530 24052 50540
rect 24108 51268 24164 51278
rect 24108 50428 24164 51212
rect 24556 51266 24612 51278
rect 24556 51214 24558 51266
rect 24610 51214 24612 51266
rect 24332 50596 24388 50606
rect 24332 50502 24388 50540
rect 23772 50372 24164 50428
rect 24444 50484 24500 50494
rect 23660 49924 23716 49934
rect 23660 49830 23716 49868
rect 23548 48974 23550 49026
rect 23602 48974 23604 49026
rect 23548 48962 23604 48974
rect 23324 48414 23326 48466
rect 23378 48414 23380 48466
rect 23324 48402 23380 48414
rect 22876 48190 22878 48242
rect 22930 48190 22932 48242
rect 22428 46674 22484 46686
rect 22428 46622 22430 46674
rect 22482 46622 22484 46674
rect 22428 45892 22484 46622
rect 22428 45826 22484 45836
rect 22260 45500 22372 45556
rect 22204 45490 22260 45500
rect 22092 44942 22094 44994
rect 22146 44942 22148 44994
rect 21868 42924 22036 42980
rect 21532 42868 21588 42878
rect 21532 42774 21588 42812
rect 21308 42754 21364 42766
rect 21308 42702 21310 42754
rect 21362 42702 21364 42754
rect 21308 42084 21364 42702
rect 21308 42018 21364 42028
rect 21532 42532 21588 42542
rect 21868 42532 21924 42542
rect 21420 41970 21476 41982
rect 21420 41918 21422 41970
rect 21474 41918 21476 41970
rect 21084 41636 21140 41646
rect 21140 41580 21364 41636
rect 21084 41570 21140 41580
rect 21196 41076 21252 41086
rect 21308 41076 21364 41580
rect 21420 41410 21476 41918
rect 21532 41970 21588 42476
rect 21644 42530 21924 42532
rect 21644 42478 21870 42530
rect 21922 42478 21924 42530
rect 21644 42476 21924 42478
rect 21644 42194 21700 42476
rect 21868 42466 21924 42476
rect 21644 42142 21646 42194
rect 21698 42142 21700 42194
rect 21644 42130 21700 42142
rect 21756 42196 21812 42206
rect 21532 41918 21534 41970
rect 21586 41918 21588 41970
rect 21532 41906 21588 41918
rect 21420 41358 21422 41410
rect 21474 41358 21476 41410
rect 21420 41346 21476 41358
rect 21756 41300 21812 42140
rect 21868 41972 21924 41982
rect 21980 41972 22036 42924
rect 22092 42644 22148 44942
rect 22316 44436 22372 44446
rect 22540 44436 22596 47068
rect 22652 47346 22708 47358
rect 22652 47294 22654 47346
rect 22706 47294 22708 47346
rect 22652 45220 22708 47294
rect 22876 46900 22932 48190
rect 23100 48132 23156 48142
rect 23156 48076 23380 48132
rect 23100 48066 23156 48076
rect 22764 46844 22932 46900
rect 22988 47460 23044 47470
rect 22764 46116 22820 46844
rect 22764 46050 22820 46060
rect 22876 46674 22932 46686
rect 22876 46622 22878 46674
rect 22930 46622 22932 46674
rect 22652 45154 22708 45164
rect 22764 45668 22820 45678
rect 22764 44996 22820 45612
rect 22316 44434 22596 44436
rect 22316 44382 22318 44434
rect 22370 44382 22596 44434
rect 22316 44380 22596 44382
rect 22652 44940 22820 44996
rect 22316 43652 22372 44380
rect 22316 43586 22372 43596
rect 22316 43428 22372 43438
rect 22316 42754 22372 43372
rect 22316 42702 22318 42754
rect 22370 42702 22372 42754
rect 22316 42690 22372 42702
rect 22092 42578 22148 42588
rect 22652 42532 22708 44940
rect 22764 43428 22820 43438
rect 22764 43334 22820 43372
rect 22876 43204 22932 46622
rect 22988 45330 23044 47404
rect 23100 47348 23156 47358
rect 23100 46002 23156 47292
rect 23212 47346 23268 47358
rect 23212 47294 23214 47346
rect 23266 47294 23268 47346
rect 23212 47124 23268 47294
rect 23212 47058 23268 47068
rect 23100 45950 23102 46002
rect 23154 45950 23156 46002
rect 23100 45938 23156 45950
rect 22988 45278 22990 45330
rect 23042 45278 23044 45330
rect 22988 45266 23044 45278
rect 22316 42476 22708 42532
rect 22764 43148 22932 43204
rect 22988 44324 23044 44334
rect 22316 42084 22372 42476
rect 22316 42018 22372 42028
rect 21868 41970 22036 41972
rect 21868 41918 21870 41970
rect 21922 41918 22036 41970
rect 21868 41916 22036 41918
rect 22428 41972 22484 41982
rect 22652 41972 22708 41982
rect 21868 41906 21924 41916
rect 22092 41858 22148 41870
rect 22092 41806 22094 41858
rect 22146 41806 22148 41858
rect 22092 41636 22148 41806
rect 22092 41570 22148 41580
rect 22316 41746 22372 41758
rect 22316 41694 22318 41746
rect 22370 41694 22372 41746
rect 22316 41412 22372 41694
rect 22316 41346 22372 41356
rect 21532 41188 21588 41198
rect 21756 41188 21812 41244
rect 21532 41186 21812 41188
rect 21532 41134 21534 41186
rect 21586 41134 21812 41186
rect 21532 41132 21812 41134
rect 22316 41188 22372 41198
rect 22428 41188 22484 41916
rect 22540 41970 22708 41972
rect 22540 41918 22654 41970
rect 22706 41918 22708 41970
rect 22540 41916 22708 41918
rect 22540 41300 22596 41916
rect 22652 41906 22708 41916
rect 22540 41206 22596 41244
rect 22652 41748 22708 41758
rect 22316 41186 22484 41188
rect 22316 41134 22318 41186
rect 22370 41134 22484 41186
rect 22316 41132 22484 41134
rect 21532 41122 21588 41132
rect 22316 41122 22372 41132
rect 21420 41076 21476 41086
rect 21308 41074 21476 41076
rect 21308 41022 21422 41074
rect 21474 41022 21476 41074
rect 21308 41020 21476 41022
rect 21196 40964 21252 41020
rect 21420 41010 21476 41020
rect 22092 41076 22148 41086
rect 21196 40908 21364 40964
rect 21196 40516 21252 40526
rect 21308 40516 21364 40908
rect 21644 40852 21700 40862
rect 21308 40460 21476 40516
rect 21196 40422 21252 40460
rect 21308 40292 21364 40302
rect 21308 39618 21364 40236
rect 21308 39566 21310 39618
rect 21362 39566 21364 39618
rect 21308 39554 21364 39566
rect 21084 39060 21140 39070
rect 21084 38164 21140 39004
rect 21084 38098 21140 38108
rect 21308 37828 21364 37838
rect 21308 37734 21364 37772
rect 21420 37380 21476 40460
rect 21644 40402 21700 40796
rect 21644 40350 21646 40402
rect 21698 40350 21700 40402
rect 21644 40338 21700 40350
rect 22092 40402 22148 41020
rect 22204 40628 22260 40638
rect 22204 40534 22260 40572
rect 22428 40626 22484 40638
rect 22428 40574 22430 40626
rect 22482 40574 22484 40626
rect 22092 40350 22094 40402
rect 22146 40350 22148 40402
rect 22092 40338 22148 40350
rect 21644 40068 21700 40078
rect 21644 39618 21700 40012
rect 22428 40068 22484 40574
rect 22652 40516 22708 41692
rect 22764 41298 22820 43148
rect 22988 43092 23044 44268
rect 23100 44100 23156 44110
rect 23100 44006 23156 44044
rect 23212 43650 23268 43662
rect 23212 43598 23214 43650
rect 23266 43598 23268 43650
rect 23212 43428 23268 43598
rect 23212 43362 23268 43372
rect 22876 43036 23044 43092
rect 23100 43314 23156 43326
rect 23100 43262 23102 43314
rect 23154 43262 23156 43314
rect 22876 41970 22932 43036
rect 22988 42754 23044 42766
rect 22988 42702 22990 42754
rect 23042 42702 23044 42754
rect 22988 42082 23044 42702
rect 22988 42030 22990 42082
rect 23042 42030 23044 42082
rect 22988 42018 23044 42030
rect 22876 41918 22878 41970
rect 22930 41918 22932 41970
rect 22876 41906 22932 41918
rect 22764 41246 22766 41298
rect 22818 41246 22820 41298
rect 22764 41234 22820 41246
rect 22876 41524 22932 41534
rect 22876 41186 22932 41468
rect 23100 41412 23156 43262
rect 23100 41346 23156 41356
rect 22876 41134 22878 41186
rect 22930 41134 22932 41186
rect 22876 41122 22932 41134
rect 23324 40740 23380 48076
rect 23772 47460 23828 50372
rect 24332 49812 24388 49822
rect 24444 49812 24500 50428
rect 24332 49810 24500 49812
rect 24332 49758 24334 49810
rect 24386 49758 24500 49810
rect 24332 49756 24500 49758
rect 24108 49364 24164 49374
rect 24108 49026 24164 49308
rect 24108 48974 24110 49026
rect 24162 48974 24164 49026
rect 24108 48962 24164 48974
rect 24220 49138 24276 49150
rect 24220 49086 24222 49138
rect 24274 49086 24276 49138
rect 24220 49028 24276 49086
rect 24220 48962 24276 48972
rect 24332 48804 24388 49756
rect 24556 49364 24612 51214
rect 24668 49924 24724 49934
rect 24668 49830 24724 49868
rect 24556 49298 24612 49308
rect 24332 48738 24388 48748
rect 24780 48580 24836 52556
rect 24892 50932 24948 54796
rect 24892 50866 24948 50876
rect 25004 50818 25060 57484
rect 26460 57204 26516 57214
rect 25564 56196 25620 56206
rect 25564 56102 25620 56140
rect 25228 55972 25284 55982
rect 25228 54514 25284 55916
rect 26124 55970 26180 55982
rect 26124 55918 26126 55970
rect 26178 55918 26180 55970
rect 26124 55412 26180 55918
rect 26124 55346 26180 55356
rect 25340 55300 25396 55310
rect 25340 54626 25396 55244
rect 26236 54740 26292 54750
rect 26236 54646 26292 54684
rect 25340 54574 25342 54626
rect 25394 54574 25396 54626
rect 25340 54562 25396 54574
rect 25228 54462 25230 54514
rect 25282 54462 25284 54514
rect 25228 53956 25284 54462
rect 26124 54514 26180 54526
rect 26124 54462 26126 54514
rect 26178 54462 26180 54514
rect 26124 54404 26180 54462
rect 26124 54338 26180 54348
rect 25228 53900 26404 53956
rect 26012 53732 26068 53742
rect 26012 53170 26068 53676
rect 26012 53118 26014 53170
rect 26066 53118 26068 53170
rect 26012 53106 26068 53118
rect 25004 50766 25006 50818
rect 25058 50766 25060 50818
rect 25004 50754 25060 50766
rect 25116 53060 25172 53070
rect 24892 50708 24948 50718
rect 24892 50614 24948 50652
rect 24332 48524 24836 48580
rect 24220 48468 24276 48478
rect 24220 48374 24276 48412
rect 23772 47366 23828 47404
rect 24108 48132 24164 48142
rect 24108 47572 24164 48076
rect 23996 46788 24052 46798
rect 23772 46676 23828 46686
rect 23772 46582 23828 46620
rect 23996 46450 24052 46732
rect 23996 46398 23998 46450
rect 24050 46398 24052 46450
rect 23996 46386 24052 46398
rect 24108 46562 24164 47516
rect 24108 46510 24110 46562
rect 24162 46510 24164 46562
rect 23884 46340 23940 46350
rect 23884 46228 23940 46284
rect 23884 46172 24052 46228
rect 23884 46004 23940 46014
rect 23884 45910 23940 45948
rect 23772 45890 23828 45902
rect 23772 45838 23774 45890
rect 23826 45838 23828 45890
rect 23660 45780 23716 45790
rect 23548 45724 23660 45780
rect 23436 45668 23492 45678
rect 23436 45574 23492 45612
rect 23436 45332 23492 45342
rect 23548 45332 23604 45724
rect 23660 45714 23716 45724
rect 23436 45330 23604 45332
rect 23436 45278 23438 45330
rect 23490 45278 23604 45330
rect 23436 45276 23604 45278
rect 23436 44548 23492 45276
rect 23436 44482 23492 44492
rect 23772 44436 23828 45838
rect 23996 45444 24052 46172
rect 24108 45778 24164 46510
rect 24108 45726 24110 45778
rect 24162 45726 24164 45778
rect 24108 45714 24164 45726
rect 23884 45332 23940 45342
rect 23996 45332 24052 45388
rect 23884 45330 24052 45332
rect 23884 45278 23886 45330
rect 23938 45278 24052 45330
rect 23884 45276 24052 45278
rect 23884 45266 23940 45276
rect 24108 45108 24164 45118
rect 23996 45106 24164 45108
rect 23996 45054 24110 45106
rect 24162 45054 24164 45106
rect 23996 45052 24164 45054
rect 23548 44100 23604 44110
rect 23548 44006 23604 44044
rect 23772 43876 23828 44380
rect 23884 44660 23940 44670
rect 23884 44322 23940 44604
rect 23996 44434 24052 45052
rect 24108 45042 24164 45052
rect 23996 44382 23998 44434
rect 24050 44382 24052 44434
rect 23996 44370 24052 44382
rect 23884 44270 23886 44322
rect 23938 44270 23940 44322
rect 23884 44258 23940 44270
rect 24108 44324 24164 44334
rect 23772 43820 23940 43876
rect 23436 43652 23492 43662
rect 23436 43558 23492 43596
rect 23772 43538 23828 43550
rect 23772 43486 23774 43538
rect 23826 43486 23828 43538
rect 23548 42756 23604 42766
rect 23436 41524 23492 41534
rect 23436 41298 23492 41468
rect 23436 41246 23438 41298
rect 23490 41246 23492 41298
rect 23436 41234 23492 41246
rect 22988 40684 23380 40740
rect 23436 40964 23492 40974
rect 22988 40626 23044 40684
rect 22988 40574 22990 40626
rect 23042 40574 23044 40626
rect 22988 40562 23044 40574
rect 22652 40450 22708 40460
rect 22428 40002 22484 40012
rect 22652 39844 22708 39854
rect 21644 39566 21646 39618
rect 21698 39566 21700 39618
rect 21644 39554 21700 39566
rect 21868 39788 22372 39844
rect 21868 38834 21924 39788
rect 22316 39732 22372 39788
rect 22428 39732 22484 39742
rect 22316 39676 22428 39732
rect 22428 39638 22484 39676
rect 21868 38782 21870 38834
rect 21922 38782 21924 38834
rect 21868 38770 21924 38782
rect 21980 39618 22036 39630
rect 21980 39566 21982 39618
rect 22034 39566 22036 39618
rect 21868 38052 21924 38062
rect 21980 38052 22036 39566
rect 22092 39620 22148 39630
rect 22092 39526 22148 39564
rect 22204 39620 22260 39630
rect 22204 39618 22372 39620
rect 22204 39566 22206 39618
rect 22258 39566 22372 39618
rect 22204 39564 22372 39566
rect 22204 39554 22260 39564
rect 22204 39396 22260 39406
rect 22204 39058 22260 39340
rect 22204 39006 22206 39058
rect 22258 39006 22260 39058
rect 22204 38994 22260 39006
rect 22316 39060 22372 39564
rect 22652 39396 22708 39788
rect 23212 39842 23268 40684
rect 23212 39790 23214 39842
rect 23266 39790 23268 39842
rect 23100 39732 23156 39742
rect 23100 39638 23156 39676
rect 22652 39330 22708 39340
rect 22428 39060 22484 39070
rect 22652 39060 22708 39070
rect 22316 39058 22708 39060
rect 22316 39006 22430 39058
rect 22482 39006 22654 39058
rect 22706 39006 22708 39058
rect 22316 39004 22708 39006
rect 22428 38994 22484 39004
rect 22652 38994 22708 39004
rect 22876 38946 22932 38958
rect 22876 38894 22878 38946
rect 22930 38894 22932 38946
rect 22316 38836 22372 38846
rect 22316 38722 22372 38780
rect 22316 38670 22318 38722
rect 22370 38670 22372 38722
rect 22316 38658 22372 38670
rect 21868 38050 22036 38052
rect 21868 37998 21870 38050
rect 21922 37998 22036 38050
rect 21868 37996 22036 37998
rect 22204 38612 22260 38622
rect 21868 37716 21924 37996
rect 21868 37650 21924 37660
rect 22092 37940 22148 37950
rect 22092 37490 22148 37884
rect 22092 37438 22094 37490
rect 22146 37438 22148 37490
rect 22092 37426 22148 37438
rect 20972 37202 21028 37212
rect 21308 37324 21476 37380
rect 21196 37042 21252 37054
rect 21196 36990 21198 37042
rect 21250 36990 21252 37042
rect 20748 36596 20804 36606
rect 20748 35028 20804 36540
rect 20748 35026 21140 35028
rect 20748 34974 20750 35026
rect 20802 34974 21140 35026
rect 20748 34972 21140 34974
rect 20748 34962 20804 34972
rect 20636 34468 20692 34748
rect 20636 34402 20692 34412
rect 20524 34188 20692 34244
rect 19852 34078 19854 34130
rect 19906 34078 19908 34130
rect 19852 34066 19908 34078
rect 19572 33740 19796 33796
rect 20188 33906 20244 33918
rect 20188 33854 20190 33906
rect 20242 33854 20244 33906
rect 19516 33730 19572 33740
rect 19516 33572 19572 33582
rect 19516 33478 19572 33516
rect 19740 33348 19796 33358
rect 20076 33348 20132 33358
rect 19628 33346 20132 33348
rect 19628 33294 19742 33346
rect 19794 33294 20078 33346
rect 20130 33294 20132 33346
rect 19628 33292 20132 33294
rect 20188 33348 20244 33854
rect 20524 33908 20580 33918
rect 20412 33348 20468 33358
rect 20188 33292 20412 33348
rect 19628 32786 19684 33292
rect 19740 33282 19796 33292
rect 20076 33282 20132 33292
rect 20412 33234 20468 33292
rect 20412 33182 20414 33234
rect 20466 33182 20468 33234
rect 20412 33170 20468 33182
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19628 32734 19630 32786
rect 19682 32734 19684 32786
rect 19628 32722 19684 32734
rect 20524 32786 20580 33852
rect 20524 32734 20526 32786
rect 20578 32734 20580 32786
rect 20524 32722 20580 32734
rect 19852 32676 19908 32686
rect 19852 32582 19908 32620
rect 19292 31666 19460 31668
rect 19292 31614 19294 31666
rect 19346 31614 19460 31666
rect 19292 31612 19460 31614
rect 19964 32562 20020 32574
rect 19964 32510 19966 32562
rect 20018 32510 20020 32562
rect 18956 30996 19012 31006
rect 18956 30902 19012 30940
rect 18620 30884 18676 30894
rect 18396 30046 18398 30098
rect 18450 30046 18452 30098
rect 18396 30034 18452 30046
rect 18508 30882 18676 30884
rect 18508 30830 18622 30882
rect 18674 30830 18676 30882
rect 18508 30828 18676 30830
rect 18508 30098 18564 30828
rect 18620 30818 18676 30828
rect 19180 30436 19236 30446
rect 19180 30210 19236 30380
rect 19180 30158 19182 30210
rect 19234 30158 19236 30210
rect 19180 30146 19236 30158
rect 18508 30046 18510 30098
rect 18562 30046 18564 30098
rect 18172 29988 18228 29998
rect 18060 29986 18228 29988
rect 18060 29934 18174 29986
rect 18226 29934 18228 29986
rect 18060 29932 18228 29934
rect 17948 29540 18004 29550
rect 17948 29446 18004 29484
rect 17836 29428 17892 29438
rect 17836 29334 17892 29372
rect 18060 29428 18116 29932
rect 18172 29922 18228 29932
rect 18060 29362 18116 29372
rect 18172 29428 18228 29438
rect 18396 29428 18452 29438
rect 18172 29426 18452 29428
rect 18172 29374 18174 29426
rect 18226 29374 18398 29426
rect 18450 29374 18452 29426
rect 18172 29372 18452 29374
rect 18172 29362 18228 29372
rect 18396 29362 18452 29372
rect 18508 29204 18564 30046
rect 19292 30100 19348 31612
rect 19964 31556 20020 32510
rect 19964 31490 20020 31500
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19404 30996 19460 31006
rect 19404 30902 19460 30940
rect 20076 30436 20132 30446
rect 19404 30212 19460 30222
rect 19404 30118 19460 30156
rect 19628 30210 19684 30222
rect 19628 30158 19630 30210
rect 19682 30158 19684 30210
rect 19292 29988 19348 30044
rect 19068 29932 19348 29988
rect 19068 29650 19124 29932
rect 19068 29598 19070 29650
rect 19122 29598 19124 29650
rect 19068 29586 19124 29598
rect 19628 29540 19684 30158
rect 20076 30212 20132 30380
rect 20076 30118 20132 30156
rect 20636 29876 20692 34188
rect 21084 34130 21140 34972
rect 21084 34078 21086 34130
rect 21138 34078 21140 34130
rect 21084 34066 21140 34078
rect 20860 33906 20916 33918
rect 20860 33854 20862 33906
rect 20914 33854 20916 33906
rect 20860 33348 20916 33854
rect 20860 33282 20916 33292
rect 21196 31892 21252 36990
rect 21308 36708 21364 37324
rect 21868 37268 21924 37278
rect 21868 37174 21924 37212
rect 21308 35700 21364 36652
rect 21420 36932 21476 36942
rect 21420 36372 21476 36876
rect 22092 36932 22148 36942
rect 22092 36706 22148 36876
rect 22092 36654 22094 36706
rect 22146 36654 22148 36706
rect 22092 36642 22148 36654
rect 21532 36596 21588 36606
rect 21532 36502 21588 36540
rect 21420 35922 21476 36316
rect 21868 36482 21924 36494
rect 21868 36430 21870 36482
rect 21922 36430 21924 36482
rect 21868 36260 21924 36430
rect 22204 36260 22260 38556
rect 22316 38164 22372 38174
rect 22316 36706 22372 38108
rect 22876 38052 22932 38894
rect 22876 37986 22932 37996
rect 22988 38834 23044 38846
rect 22988 38782 22990 38834
rect 23042 38782 23044 38834
rect 22988 37940 23044 38782
rect 22988 37604 23044 37884
rect 22988 37538 23044 37548
rect 22316 36654 22318 36706
rect 22370 36654 22372 36706
rect 22316 36596 22372 36654
rect 22316 36530 22372 36540
rect 22876 36484 22932 36494
rect 22764 36482 22932 36484
rect 22764 36430 22878 36482
rect 22930 36430 22932 36482
rect 22764 36428 22932 36430
rect 22764 36370 22820 36428
rect 22876 36418 22932 36428
rect 22764 36318 22766 36370
rect 22818 36318 22820 36370
rect 22764 36306 22820 36318
rect 21868 36204 22260 36260
rect 21420 35870 21422 35922
rect 21474 35870 21476 35922
rect 21420 35858 21476 35870
rect 21308 35634 21364 35644
rect 22092 35140 22148 36204
rect 22764 35812 22820 35822
rect 22764 35718 22820 35756
rect 23212 35308 23268 39790
rect 23324 40068 23380 40078
rect 23324 39284 23380 40012
rect 23436 39842 23492 40908
rect 23436 39790 23438 39842
rect 23490 39790 23492 39842
rect 23436 39778 23492 39790
rect 23324 39218 23380 39228
rect 23548 38668 23604 42700
rect 23660 42084 23716 42094
rect 23660 41990 23716 42028
rect 23772 40402 23828 43486
rect 23884 43540 23940 43820
rect 23884 43474 23940 43484
rect 23884 43204 23940 43214
rect 23884 42756 23940 43148
rect 24108 43204 24164 44268
rect 24332 43652 24388 48524
rect 24668 48356 24724 48366
rect 24556 48300 24668 48356
rect 24444 45780 24500 45790
rect 24444 45686 24500 45724
rect 24444 45220 24500 45230
rect 24444 45126 24500 45164
rect 24556 44548 24612 48300
rect 24668 48262 24724 48300
rect 24668 47572 24724 47582
rect 24668 47478 24724 47516
rect 25116 47460 25172 53004
rect 25564 52836 25620 52846
rect 25340 52780 25564 52836
rect 25228 51604 25284 51614
rect 25228 51510 25284 51548
rect 25228 51380 25284 51390
rect 25228 48132 25284 51324
rect 25340 49812 25396 52780
rect 25564 52742 25620 52780
rect 26012 52388 26068 52398
rect 25676 52164 25732 52174
rect 25676 51490 25732 52108
rect 26012 52162 26068 52332
rect 26012 52110 26014 52162
rect 26066 52110 26068 52162
rect 26012 52098 26068 52110
rect 25676 51438 25678 51490
rect 25730 51438 25732 51490
rect 25452 51378 25508 51390
rect 25452 51326 25454 51378
rect 25506 51326 25508 51378
rect 25452 50428 25508 51326
rect 25564 51154 25620 51166
rect 25564 51102 25566 51154
rect 25618 51102 25620 51154
rect 25564 50596 25620 51102
rect 25564 50530 25620 50540
rect 25452 50372 25620 50428
rect 25564 49924 25620 50372
rect 25676 50148 25732 51438
rect 26124 52052 26180 52062
rect 26124 51380 26180 51996
rect 26124 51286 26180 51324
rect 26124 50820 26180 50830
rect 25788 50708 25844 50718
rect 25788 50260 25844 50652
rect 25900 50260 25956 50270
rect 25788 50204 25900 50260
rect 25900 50194 25956 50204
rect 25676 50082 25732 50092
rect 26012 50148 26068 50158
rect 25452 49812 25508 49822
rect 25340 49810 25508 49812
rect 25340 49758 25454 49810
rect 25506 49758 25508 49810
rect 25340 49756 25508 49758
rect 25452 48692 25508 49756
rect 25564 48916 25620 49868
rect 26012 49476 26068 50092
rect 26012 49028 26068 49420
rect 26012 48962 26068 48972
rect 25676 48916 25732 48926
rect 25564 48860 25676 48916
rect 25676 48850 25732 48860
rect 25900 48804 25956 48814
rect 25452 48636 25732 48692
rect 25564 48244 25620 48254
rect 25452 48132 25508 48142
rect 25228 48130 25508 48132
rect 25228 48078 25454 48130
rect 25506 48078 25508 48130
rect 25228 48076 25508 48078
rect 25340 47908 25396 47918
rect 24780 47458 25172 47460
rect 24780 47406 25118 47458
rect 25170 47406 25172 47458
rect 24780 47404 25172 47406
rect 24780 47348 24836 47404
rect 25116 47394 25172 47404
rect 25228 47460 25284 47470
rect 24668 47292 24836 47348
rect 24668 46340 24724 47292
rect 25228 47236 25284 47404
rect 25340 47458 25396 47852
rect 25340 47406 25342 47458
rect 25394 47406 25396 47458
rect 25340 47394 25396 47406
rect 25452 47348 25508 48076
rect 25564 47570 25620 48188
rect 25676 47908 25732 48636
rect 25788 48242 25844 48254
rect 25788 48190 25790 48242
rect 25842 48190 25844 48242
rect 25788 48020 25844 48190
rect 25788 47954 25844 47964
rect 25676 47842 25732 47852
rect 25564 47518 25566 47570
rect 25618 47518 25620 47570
rect 25564 47506 25620 47518
rect 25676 47684 25732 47694
rect 25452 47282 25508 47292
rect 25676 47346 25732 47628
rect 25676 47294 25678 47346
rect 25730 47294 25732 47346
rect 25228 47180 25396 47236
rect 24668 45890 24724 46284
rect 24892 46676 24948 46686
rect 24780 46116 24836 46126
rect 24780 46002 24836 46060
rect 24780 45950 24782 46002
rect 24834 45950 24836 46002
rect 24780 45938 24836 45950
rect 24668 45838 24670 45890
rect 24722 45838 24724 45890
rect 24668 45826 24724 45838
rect 24668 45444 24724 45454
rect 24668 45330 24724 45388
rect 24668 45278 24670 45330
rect 24722 45278 24724 45330
rect 24668 45266 24724 45278
rect 24780 45220 24836 45230
rect 24780 45126 24836 45164
rect 24556 44482 24612 44492
rect 24892 44546 24948 46620
rect 25228 46562 25284 46574
rect 25228 46510 25230 46562
rect 25282 46510 25284 46562
rect 25228 46116 25284 46510
rect 25228 46050 25284 46060
rect 25116 45666 25172 45678
rect 25116 45614 25118 45666
rect 25170 45614 25172 45666
rect 25116 45108 25172 45614
rect 25340 45668 25396 47180
rect 25676 46788 25732 47294
rect 25900 46900 25956 48748
rect 26124 48354 26180 50764
rect 26236 50372 26292 50382
rect 26236 49026 26292 50316
rect 26236 48974 26238 49026
rect 26290 48974 26292 49026
rect 26236 48962 26292 48974
rect 26124 48302 26126 48354
rect 26178 48302 26180 48354
rect 26012 47460 26068 47498
rect 26012 47394 26068 47404
rect 25900 46844 26068 46900
rect 25676 46732 25956 46788
rect 25564 46564 25620 46574
rect 25340 45602 25396 45612
rect 25452 46450 25508 46462
rect 25452 46398 25454 46450
rect 25506 46398 25508 46450
rect 25340 45444 25396 45454
rect 25340 45330 25396 45388
rect 25340 45278 25342 45330
rect 25394 45278 25396 45330
rect 25340 45266 25396 45278
rect 25452 45220 25508 46398
rect 25452 45154 25508 45164
rect 25116 45042 25172 45052
rect 24892 44494 24894 44546
rect 24946 44494 24948 44546
rect 24892 44436 24948 44494
rect 24892 44370 24948 44380
rect 25228 44660 25284 44670
rect 24332 43558 24388 43596
rect 24556 44324 24612 44334
rect 24108 43138 24164 43148
rect 23884 42690 23940 42700
rect 24444 42756 24500 42766
rect 24444 42662 24500 42700
rect 24108 42530 24164 42542
rect 24108 42478 24110 42530
rect 24162 42478 24164 42530
rect 24108 42420 24164 42478
rect 24108 42354 24164 42364
rect 23772 40350 23774 40402
rect 23826 40350 23828 40402
rect 23436 38612 23604 38668
rect 23660 39618 23716 39630
rect 23660 39566 23662 39618
rect 23714 39566 23716 39618
rect 23660 38668 23716 39566
rect 23772 38948 23828 40350
rect 23772 38882 23828 38892
rect 23884 41970 23940 41982
rect 23884 41918 23886 41970
rect 23938 41918 23940 41970
rect 23884 38724 23940 41918
rect 24220 41636 24276 41646
rect 24220 41298 24276 41580
rect 24220 41246 24222 41298
rect 24274 41246 24276 41298
rect 24220 41234 24276 41246
rect 24556 41188 24612 44268
rect 25004 44324 25060 44334
rect 25004 44230 25060 44268
rect 24892 43652 24948 43662
rect 24892 42642 24948 43596
rect 24892 42590 24894 42642
rect 24946 42590 24948 42642
rect 24892 42578 24948 42590
rect 24332 41186 24612 41188
rect 24332 41134 24558 41186
rect 24610 41134 24612 41186
rect 24332 41132 24612 41134
rect 24220 41076 24276 41086
rect 24220 39732 24276 41020
rect 24332 40404 24388 41132
rect 24556 41122 24612 41132
rect 25228 41972 25284 44604
rect 25340 44210 25396 44222
rect 25340 44158 25342 44210
rect 25394 44158 25396 44210
rect 25340 44100 25396 44158
rect 25340 44034 25396 44044
rect 25564 43764 25620 46508
rect 25788 46450 25844 46462
rect 25788 46398 25790 46450
rect 25842 46398 25844 46450
rect 25788 46228 25844 46398
rect 25788 46162 25844 46172
rect 25676 45890 25732 45902
rect 25676 45838 25678 45890
rect 25730 45838 25732 45890
rect 25676 45780 25732 45838
rect 25676 45714 25732 45724
rect 25900 45556 25956 46732
rect 25452 43708 25620 43764
rect 25676 45500 25956 45556
rect 25340 43540 25396 43550
rect 25340 43446 25396 43484
rect 25340 41972 25396 41982
rect 25228 41970 25396 41972
rect 25228 41918 25342 41970
rect 25394 41918 25396 41970
rect 25228 41916 25396 41918
rect 24780 40964 24836 40974
rect 24780 40870 24836 40908
rect 24332 40310 24388 40348
rect 25004 40180 25060 40190
rect 24220 39730 24500 39732
rect 24220 39678 24222 39730
rect 24274 39678 24500 39730
rect 24220 39676 24500 39678
rect 24220 39666 24276 39676
rect 24444 39620 24500 39676
rect 25004 39730 25060 40124
rect 25004 39678 25006 39730
rect 25058 39678 25060 39730
rect 25004 39666 25060 39678
rect 24444 39618 24612 39620
rect 24444 39566 24446 39618
rect 24498 39566 24612 39618
rect 24444 39564 24612 39566
rect 24444 39554 24500 39564
rect 23996 39396 24052 39406
rect 23996 39058 24052 39340
rect 24220 39172 24276 39182
rect 23996 39006 23998 39058
rect 24050 39006 24052 39058
rect 23996 38994 24052 39006
rect 24108 39060 24164 39070
rect 24108 38834 24164 39004
rect 24108 38782 24110 38834
rect 24162 38782 24164 38834
rect 24108 38770 24164 38782
rect 23660 38612 23828 38668
rect 23884 38658 23940 38668
rect 23996 38722 24052 38734
rect 23996 38670 23998 38722
rect 24050 38670 24052 38722
rect 23436 38052 23492 38612
rect 23436 37958 23492 37996
rect 23548 37828 23604 37838
rect 23548 37490 23604 37772
rect 23548 37438 23550 37490
rect 23602 37438 23604 37490
rect 23548 37380 23604 37438
rect 23548 37314 23604 37324
rect 23548 36594 23604 36606
rect 23548 36542 23550 36594
rect 23602 36542 23604 36594
rect 23100 35252 23268 35308
rect 23324 36036 23380 36046
rect 22428 35140 22484 35150
rect 22092 35084 22428 35140
rect 21980 35028 22036 35038
rect 21868 34972 21980 35028
rect 21308 34916 21364 34926
rect 21308 34130 21364 34860
rect 21868 34914 21924 34972
rect 21980 34962 22036 34972
rect 22316 35026 22372 35084
rect 22428 35074 22484 35084
rect 22316 34974 22318 35026
rect 22370 34974 22372 35026
rect 22316 34962 22372 34974
rect 22764 35028 22820 35038
rect 22764 34916 22820 34972
rect 21868 34862 21870 34914
rect 21922 34862 21924 34914
rect 21868 34850 21924 34862
rect 22428 34914 22820 34916
rect 22428 34862 22766 34914
rect 22818 34862 22820 34914
rect 22428 34860 22820 34862
rect 21532 34692 21588 34702
rect 21308 34078 21310 34130
rect 21362 34078 21364 34130
rect 21308 33908 21364 34078
rect 21308 33842 21364 33852
rect 21420 34356 21476 34366
rect 21532 34356 21588 34636
rect 21644 34356 21700 34366
rect 21532 34354 21700 34356
rect 21532 34302 21646 34354
rect 21698 34302 21700 34354
rect 21532 34300 21700 34302
rect 21420 33460 21476 34300
rect 21644 34290 21700 34300
rect 21756 34356 21812 34366
rect 21756 34262 21812 34300
rect 22428 34354 22484 34860
rect 22764 34850 22820 34860
rect 22428 34302 22430 34354
rect 22482 34302 22484 34354
rect 22428 34290 22484 34302
rect 22988 34690 23044 34702
rect 22988 34638 22990 34690
rect 23042 34638 23044 34690
rect 22988 34356 23044 34638
rect 22988 34290 23044 34300
rect 21532 34132 21588 34142
rect 21532 34038 21588 34076
rect 21532 33460 21588 33470
rect 21420 33458 21588 33460
rect 21420 33406 21534 33458
rect 21586 33406 21588 33458
rect 21420 33404 21588 33406
rect 21532 33394 21588 33404
rect 22988 33460 23044 33470
rect 23100 33460 23156 35252
rect 23212 34356 23268 34366
rect 23324 34356 23380 35980
rect 23548 35924 23604 36542
rect 23548 35858 23604 35868
rect 23548 34468 23604 34478
rect 23212 34354 23492 34356
rect 23212 34302 23214 34354
rect 23266 34302 23492 34354
rect 23212 34300 23492 34302
rect 23212 34290 23268 34300
rect 22988 33458 23156 33460
rect 22988 33406 22990 33458
rect 23042 33406 23156 33458
rect 22988 33404 23156 33406
rect 23436 33572 23492 34300
rect 23548 34354 23604 34412
rect 23548 34302 23550 34354
rect 23602 34302 23604 34354
rect 23548 34290 23604 34302
rect 23660 34356 23716 34366
rect 23772 34356 23828 38556
rect 23996 38164 24052 38670
rect 24220 38668 24276 39116
rect 23884 38108 24052 38164
rect 24108 38612 24276 38668
rect 23884 36148 23940 38108
rect 23996 37940 24052 37950
rect 24108 37940 24164 38612
rect 24556 38164 24612 39564
rect 25116 39508 25172 39518
rect 25116 39414 25172 39452
rect 24892 39394 24948 39406
rect 24892 39342 24894 39394
rect 24946 39342 24948 39394
rect 24892 38612 24948 39342
rect 25228 38668 25284 41916
rect 25340 41906 25396 41916
rect 25452 41412 25508 43708
rect 25564 43538 25620 43550
rect 25564 43486 25566 43538
rect 25618 43486 25620 43538
rect 25564 43092 25620 43486
rect 25564 43026 25620 43036
rect 25676 42756 25732 45500
rect 25788 45332 25844 45342
rect 26012 45332 26068 46844
rect 25788 45330 26068 45332
rect 25788 45278 25790 45330
rect 25842 45278 26068 45330
rect 25788 45276 26068 45278
rect 25788 43652 25844 45276
rect 25788 43586 25844 43596
rect 26124 43652 26180 48302
rect 26348 47572 26404 53900
rect 26460 53730 26516 57148
rect 26684 57204 26740 57820
rect 30604 57652 30660 57662
rect 26684 57138 26740 57148
rect 27580 57316 27636 57326
rect 27020 56644 27076 56654
rect 27020 56306 27076 56588
rect 27020 56254 27022 56306
rect 27074 56254 27076 56306
rect 27020 56242 27076 56254
rect 26796 55970 26852 55982
rect 26796 55918 26798 55970
rect 26850 55918 26852 55970
rect 26796 55636 26852 55918
rect 27580 55970 27636 57260
rect 27580 55918 27582 55970
rect 27634 55918 27636 55970
rect 26796 55580 26964 55636
rect 26684 55412 26740 55422
rect 26684 55298 26740 55356
rect 26684 55246 26686 55298
rect 26738 55246 26740 55298
rect 26684 55234 26740 55246
rect 26796 55410 26852 55422
rect 26796 55358 26798 55410
rect 26850 55358 26852 55410
rect 26796 54852 26852 55358
rect 26908 55300 26964 55580
rect 27580 55300 27636 55918
rect 28476 56194 28532 56206
rect 28476 56142 28478 56194
rect 28530 56142 28532 56194
rect 28364 55860 28420 55870
rect 26908 55244 27076 55300
rect 26796 54786 26852 54796
rect 26908 54516 26964 54526
rect 26908 54422 26964 54460
rect 26460 53678 26462 53730
rect 26514 53678 26516 53730
rect 26460 53620 26516 53678
rect 26460 53554 26516 53564
rect 26684 53732 26740 53742
rect 26572 53508 26628 53518
rect 26572 53396 26628 53452
rect 26460 53340 26628 53396
rect 26460 52500 26516 53340
rect 26572 52836 26628 52846
rect 26572 52742 26628 52780
rect 26460 51044 26516 52444
rect 26684 52388 26740 53676
rect 26908 53508 26964 53518
rect 27020 53508 27076 55244
rect 27580 55234 27636 55244
rect 27692 55858 28420 55860
rect 27692 55806 28366 55858
rect 28418 55806 28420 55858
rect 27692 55804 28420 55806
rect 27580 55076 27636 55086
rect 27580 54180 27636 55020
rect 27580 54114 27636 54124
rect 27692 53730 27748 55804
rect 28364 55794 28420 55804
rect 27692 53678 27694 53730
rect 27746 53678 27748 53730
rect 27692 53666 27748 53678
rect 27916 55636 27972 55646
rect 27916 55186 27972 55580
rect 28364 55524 28420 55534
rect 28476 55524 28532 56142
rect 28700 56196 28756 56206
rect 28700 55860 28756 56140
rect 28700 55794 28756 55804
rect 29596 55970 29652 55982
rect 29596 55918 29598 55970
rect 29650 55918 29652 55970
rect 28420 55468 28532 55524
rect 29484 55748 29540 55758
rect 28364 55458 28420 55468
rect 27916 55134 27918 55186
rect 27970 55134 27972 55186
rect 26964 53452 27076 53508
rect 27356 53506 27412 53518
rect 27356 53454 27358 53506
rect 27410 53454 27412 53506
rect 26908 53442 26964 53452
rect 27356 52948 27412 53454
rect 27916 53284 27972 55134
rect 28252 55300 28308 55310
rect 28140 54514 28196 54526
rect 28140 54462 28142 54514
rect 28194 54462 28196 54514
rect 28140 54068 28196 54462
rect 28140 53844 28196 54012
rect 28140 53778 28196 53788
rect 28028 53508 28084 53518
rect 28028 53414 28084 53452
rect 28252 53396 28308 55244
rect 28476 55186 28532 55198
rect 28476 55134 28478 55186
rect 28530 55134 28532 55186
rect 28364 55074 28420 55086
rect 28364 55022 28366 55074
rect 28418 55022 28420 55074
rect 28364 54516 28420 55022
rect 28364 54450 28420 54460
rect 28140 53340 28308 53396
rect 28364 54292 28420 54302
rect 28364 53730 28420 54236
rect 28364 53678 28366 53730
rect 28418 53678 28420 53730
rect 28364 53396 28420 53678
rect 27916 53228 28084 53284
rect 28028 53172 28084 53228
rect 28028 53106 28084 53116
rect 27916 53058 27972 53070
rect 27916 53006 27918 53058
rect 27970 53006 27972 53058
rect 27412 52892 27524 52948
rect 27356 52882 27412 52892
rect 26684 52322 26740 52332
rect 27020 52834 27076 52846
rect 27020 52782 27022 52834
rect 27074 52782 27076 52834
rect 26796 52276 26852 52286
rect 26852 52220 26964 52276
rect 26796 52210 26852 52220
rect 26908 51490 26964 52220
rect 26908 51438 26910 51490
rect 26962 51438 26964 51490
rect 26908 51426 26964 51438
rect 26572 51268 26628 51278
rect 26572 51174 26628 51212
rect 27020 51156 27076 52782
rect 27132 52164 27188 52174
rect 27132 52070 27188 52108
rect 27132 51380 27188 51390
rect 27132 51286 27188 51324
rect 26908 51100 27076 51156
rect 26460 50988 26740 51044
rect 26460 50482 26516 50494
rect 26460 50430 26462 50482
rect 26514 50430 26516 50482
rect 26460 50148 26516 50430
rect 26460 50082 26516 50092
rect 26572 49924 26628 49934
rect 26236 47516 26404 47572
rect 26460 49868 26572 49924
rect 26236 47124 26292 47516
rect 26348 47348 26404 47358
rect 26348 47254 26404 47292
rect 26236 47012 26404 47124
rect 26236 46676 26292 47012
rect 26236 46610 26292 46620
rect 26460 46676 26516 49868
rect 26572 49830 26628 49868
rect 26572 49028 26628 49038
rect 26572 48468 26628 48972
rect 26684 48804 26740 50988
rect 26908 50596 26964 51100
rect 27468 50820 27524 52892
rect 27580 52612 27636 52622
rect 27580 52274 27636 52556
rect 27580 52222 27582 52274
rect 27634 52222 27636 52274
rect 27580 52210 27636 52222
rect 27916 52276 27972 53006
rect 28028 52500 28084 52510
rect 28028 52386 28084 52444
rect 28028 52334 28030 52386
rect 28082 52334 28084 52386
rect 28028 52322 28084 52334
rect 27916 52210 27972 52220
rect 27244 50764 27524 50820
rect 27804 51268 27860 51278
rect 26908 50540 27076 50596
rect 26796 50372 26852 50382
rect 26796 49812 26852 50316
rect 26908 50370 26964 50382
rect 26908 50318 26910 50370
rect 26962 50318 26964 50370
rect 26908 50148 26964 50318
rect 26908 50082 26964 50092
rect 26796 49746 26852 49756
rect 26796 49588 26852 49598
rect 26796 49138 26852 49532
rect 26796 49086 26798 49138
rect 26850 49086 26852 49138
rect 26796 49074 26852 49086
rect 26908 49364 26964 49374
rect 26684 48738 26740 48748
rect 26796 48468 26852 48506
rect 26628 48412 26740 48468
rect 26572 48402 26628 48412
rect 26572 48020 26628 48030
rect 26572 47346 26628 47964
rect 26572 47294 26574 47346
rect 26626 47294 26628 47346
rect 26572 47282 26628 47294
rect 26460 46610 26516 46620
rect 26684 46676 26740 48412
rect 26796 48402 26852 48412
rect 26796 48242 26852 48254
rect 26796 48190 26798 48242
rect 26850 48190 26852 48242
rect 26796 47908 26852 48190
rect 26796 47842 26852 47852
rect 26684 46610 26740 46620
rect 26572 46564 26628 46574
rect 26572 46470 26628 46508
rect 26236 46452 26292 46462
rect 26236 46002 26292 46396
rect 26796 46452 26852 46462
rect 26796 46004 26852 46396
rect 26236 45950 26238 46002
rect 26290 45950 26292 46002
rect 26236 45938 26292 45950
rect 26684 45948 26852 46004
rect 26572 45892 26628 45930
rect 26572 45826 26628 45836
rect 26572 45444 26628 45454
rect 26236 44996 26292 45006
rect 26236 44902 26292 44940
rect 26460 44322 26516 44334
rect 26460 44270 26462 44322
rect 26514 44270 26516 44322
rect 26460 44212 26516 44270
rect 26460 44146 26516 44156
rect 26572 44100 26628 45388
rect 26684 45108 26740 45948
rect 26908 45444 26964 49308
rect 27020 49028 27076 50540
rect 27244 50428 27300 50764
rect 27356 50596 27412 50606
rect 27356 50502 27412 50540
rect 27132 50372 27300 50428
rect 27468 50482 27524 50494
rect 27468 50430 27470 50482
rect 27522 50430 27524 50482
rect 27356 50372 27412 50382
rect 27132 50306 27188 50316
rect 27244 50148 27300 50158
rect 27356 50148 27412 50316
rect 27300 50092 27412 50148
rect 27468 50148 27524 50430
rect 27244 50082 27300 50092
rect 27468 50082 27524 50092
rect 27244 49812 27300 49822
rect 27244 49718 27300 49756
rect 27804 49810 27860 51212
rect 27804 49758 27806 49810
rect 27858 49758 27860 49810
rect 27804 49700 27860 49758
rect 27804 49634 27860 49644
rect 27916 50820 27972 50830
rect 27244 49028 27300 49038
rect 27020 49026 27300 49028
rect 27020 48974 27246 49026
rect 27298 48974 27300 49026
rect 27020 48972 27300 48974
rect 27244 48468 27300 48972
rect 27804 49028 27860 49038
rect 27916 49028 27972 50764
rect 28028 50594 28084 50606
rect 28028 50542 28030 50594
rect 28082 50542 28084 50594
rect 28028 49812 28084 50542
rect 28028 49746 28084 49756
rect 28028 49028 28084 49038
rect 27916 49026 28084 49028
rect 27916 48974 28030 49026
rect 28082 48974 28084 49026
rect 27916 48972 28084 48974
rect 27356 48916 27412 48926
rect 27356 48822 27412 48860
rect 27580 48802 27636 48814
rect 27580 48750 27582 48802
rect 27634 48750 27636 48802
rect 27468 48468 27524 48478
rect 27244 48466 27524 48468
rect 27244 48414 27470 48466
rect 27522 48414 27524 48466
rect 27244 48412 27524 48414
rect 27468 48356 27524 48412
rect 27244 48244 27300 48254
rect 27244 48150 27300 48188
rect 27244 47572 27300 47582
rect 27244 47478 27300 47516
rect 27468 47012 27524 48300
rect 27580 48354 27636 48750
rect 27580 48302 27582 48354
rect 27634 48302 27636 48354
rect 27580 48290 27636 48302
rect 27692 48802 27748 48814
rect 27692 48750 27694 48802
rect 27746 48750 27748 48802
rect 27692 48354 27748 48750
rect 27804 48804 27860 48972
rect 28028 48962 28084 48972
rect 27916 48804 27972 48814
rect 27804 48802 27972 48804
rect 27804 48750 27918 48802
rect 27970 48750 27972 48802
rect 27804 48748 27972 48750
rect 27916 48738 27972 48748
rect 28028 48804 28084 48814
rect 28028 48580 28084 48748
rect 27692 48302 27694 48354
rect 27746 48302 27748 48354
rect 27692 48244 27748 48302
rect 27692 48178 27748 48188
rect 27804 48524 28084 48580
rect 27468 46946 27524 46956
rect 27580 48020 27636 48030
rect 27468 46788 27524 46798
rect 27468 46694 27524 46732
rect 27020 46562 27076 46574
rect 27020 46510 27022 46562
rect 27074 46510 27076 46562
rect 27020 46452 27076 46510
rect 27020 46386 27076 46396
rect 27468 46452 27524 46462
rect 27356 46004 27412 46014
rect 27244 46002 27412 46004
rect 27244 45950 27358 46002
rect 27410 45950 27412 46002
rect 27244 45948 27412 45950
rect 27020 45780 27076 45790
rect 27020 45686 27076 45724
rect 26908 45378 26964 45388
rect 27020 45108 27076 45118
rect 27244 45108 27300 45948
rect 27356 45938 27412 45948
rect 27356 45778 27412 45790
rect 27356 45726 27358 45778
rect 27410 45726 27412 45778
rect 27356 45668 27412 45726
rect 27356 45602 27412 45612
rect 26684 45106 26964 45108
rect 26684 45054 26686 45106
rect 26738 45054 26964 45106
rect 26684 45052 26964 45054
rect 26684 45042 26740 45052
rect 26796 44324 26852 44334
rect 26796 44230 26852 44268
rect 26572 44044 26852 44100
rect 26124 43586 26180 43596
rect 26572 43538 26628 43550
rect 26572 43486 26574 43538
rect 26626 43486 26628 43538
rect 26348 43428 26404 43438
rect 25900 43204 25956 43214
rect 25676 42700 25844 42756
rect 25340 41356 25508 41412
rect 25564 42084 25620 42094
rect 25340 40852 25396 41356
rect 25340 40786 25396 40796
rect 25452 41186 25508 41198
rect 25452 41134 25454 41186
rect 25506 41134 25508 41186
rect 25340 40402 25396 40414
rect 25340 40350 25342 40402
rect 25394 40350 25396 40402
rect 25340 39508 25396 40350
rect 25452 39620 25508 41134
rect 25564 41076 25620 42028
rect 25676 41860 25732 41870
rect 25676 41766 25732 41804
rect 25564 41010 25620 41020
rect 25676 40964 25732 40974
rect 25676 40870 25732 40908
rect 25788 40740 25844 42700
rect 25900 42754 25956 43148
rect 26348 42868 26404 43372
rect 26348 42802 26404 42812
rect 26460 43314 26516 43326
rect 26460 43262 26462 43314
rect 26514 43262 26516 43314
rect 25900 42702 25902 42754
rect 25954 42702 25956 42754
rect 25900 42690 25956 42702
rect 26012 42642 26068 42654
rect 26012 42590 26014 42642
rect 26066 42590 26068 42642
rect 25900 42084 25956 42094
rect 26012 42084 26068 42590
rect 25956 42028 26068 42084
rect 26348 42308 26404 42318
rect 25900 42018 25956 42028
rect 26012 41412 26068 41422
rect 26012 41318 26068 41356
rect 26348 41412 26404 42252
rect 26460 42196 26516 43262
rect 26572 42868 26628 43486
rect 26572 42774 26628 42812
rect 26796 43540 26852 44044
rect 26796 42754 26852 43484
rect 26796 42702 26798 42754
rect 26850 42702 26852 42754
rect 26796 42690 26852 42702
rect 26908 42308 26964 45052
rect 27020 45106 27300 45108
rect 27020 45054 27022 45106
rect 27074 45054 27300 45106
rect 27020 45052 27300 45054
rect 27356 45444 27412 45454
rect 27020 44100 27076 45052
rect 27020 44034 27076 44044
rect 27020 43652 27076 43662
rect 27020 43558 27076 43596
rect 26908 42242 26964 42252
rect 26796 42196 26852 42206
rect 26460 42140 26628 42196
rect 26460 41970 26516 41982
rect 26460 41918 26462 41970
rect 26514 41918 26516 41970
rect 26460 41636 26516 41918
rect 26572 41748 26628 42140
rect 26572 41682 26628 41692
rect 27356 42196 27412 45388
rect 27468 44884 27524 46396
rect 27468 44818 27524 44828
rect 27580 44660 27636 47964
rect 27692 47684 27748 47694
rect 27692 47570 27748 47628
rect 27692 47518 27694 47570
rect 27746 47518 27748 47570
rect 27692 47506 27748 47518
rect 27692 46900 27748 46910
rect 27692 45890 27748 46844
rect 27692 45838 27694 45890
rect 27746 45838 27748 45890
rect 27692 45444 27748 45838
rect 27692 45378 27748 45388
rect 27468 44604 27636 44660
rect 27804 45218 27860 48524
rect 28028 48356 28084 48366
rect 28028 48130 28084 48300
rect 28028 48078 28030 48130
rect 28082 48078 28084 48130
rect 28028 48066 28084 48078
rect 28028 47348 28084 47358
rect 28028 47254 28084 47292
rect 27916 47124 27972 47134
rect 27916 46674 27972 47068
rect 27916 46622 27918 46674
rect 27970 46622 27972 46674
rect 27916 46610 27972 46622
rect 28028 46004 28084 46014
rect 27804 45166 27806 45218
rect 27858 45166 27860 45218
rect 27468 43092 27524 44604
rect 27804 44212 27860 45166
rect 27916 45948 28028 46004
rect 27916 45106 27972 45948
rect 28028 45938 28084 45948
rect 27916 45054 27918 45106
rect 27970 45054 27972 45106
rect 27916 45042 27972 45054
rect 28028 44996 28084 45006
rect 28028 44902 28084 44940
rect 27804 44146 27860 44156
rect 27468 43026 27524 43036
rect 27580 43652 27636 43662
rect 27468 42868 27524 42878
rect 27468 42774 27524 42812
rect 27580 42756 27636 43596
rect 28028 43540 28084 43550
rect 28140 43540 28196 53340
rect 28364 53330 28420 53340
rect 28476 52946 28532 55134
rect 29260 55076 29316 55086
rect 29260 54982 29316 55020
rect 29484 54514 29540 55692
rect 29484 54462 29486 54514
rect 29538 54462 29540 54514
rect 29484 54450 29540 54462
rect 29596 53956 29652 55918
rect 30156 55970 30212 55982
rect 30156 55918 30158 55970
rect 30210 55918 30212 55970
rect 29820 55298 29876 55310
rect 29820 55246 29822 55298
rect 29874 55246 29876 55298
rect 29820 55076 29876 55246
rect 29596 53890 29652 53900
rect 29708 54402 29764 54414
rect 29708 54350 29710 54402
rect 29762 54350 29764 54402
rect 28476 52894 28478 52946
rect 28530 52894 28532 52946
rect 28252 52612 28308 52622
rect 28252 49812 28308 52556
rect 28476 52500 28532 52894
rect 28588 53618 28644 53630
rect 28588 53566 28590 53618
rect 28642 53566 28644 53618
rect 28588 52612 28644 53566
rect 29148 53620 29204 53630
rect 29148 53526 29204 53564
rect 29596 53620 29652 53630
rect 29484 53508 29540 53518
rect 29372 53506 29540 53508
rect 29372 53454 29486 53506
rect 29538 53454 29540 53506
rect 29372 53452 29540 53454
rect 29036 53060 29092 53070
rect 28924 52836 28980 52846
rect 28924 52742 28980 52780
rect 28588 52546 28644 52556
rect 28476 52434 28532 52444
rect 29036 52162 29092 53004
rect 29036 52110 29038 52162
rect 29090 52110 29092 52162
rect 29036 52098 29092 52110
rect 29372 51940 29428 53452
rect 29484 53442 29540 53452
rect 29484 53172 29540 53182
rect 29484 52946 29540 53116
rect 29484 52894 29486 52946
rect 29538 52894 29540 52946
rect 29484 52882 29540 52894
rect 29596 52274 29652 53564
rect 29596 52222 29598 52274
rect 29650 52222 29652 52274
rect 29596 52210 29652 52222
rect 29708 52164 29764 54350
rect 29820 53618 29876 55020
rect 30156 54404 30212 55918
rect 30156 54338 30212 54348
rect 30268 55410 30324 55422
rect 30268 55358 30270 55410
rect 30322 55358 30324 55410
rect 30268 54292 30324 55358
rect 30380 54628 30436 54638
rect 30436 54572 30548 54628
rect 30380 54562 30436 54572
rect 30268 54226 30324 54236
rect 30380 54180 30436 54190
rect 29820 53566 29822 53618
rect 29874 53566 29876 53618
rect 29820 53396 29876 53566
rect 29932 53956 29988 53966
rect 29932 53618 29988 53900
rect 30156 53732 30212 53742
rect 30156 53638 30212 53676
rect 29932 53566 29934 53618
rect 29986 53566 29988 53618
rect 29932 53554 29988 53566
rect 29820 53330 29876 53340
rect 30380 52948 30436 54124
rect 30492 53060 30548 54572
rect 30604 54292 30660 57596
rect 30716 56084 30772 56094
rect 30716 55990 30772 56028
rect 30940 55972 30996 59200
rect 36316 57764 36372 57774
rect 34300 56308 34356 56318
rect 34356 56252 34468 56308
rect 34300 56242 34356 56252
rect 31500 56082 31556 56094
rect 31500 56030 31502 56082
rect 31554 56030 31556 56082
rect 30940 55906 30996 55916
rect 31052 55970 31108 55982
rect 31052 55918 31054 55970
rect 31106 55918 31108 55970
rect 31052 55188 31108 55918
rect 31052 55122 31108 55132
rect 31164 55300 31220 55310
rect 31500 55300 31556 56030
rect 34300 56082 34356 56094
rect 34300 56030 34302 56082
rect 34354 56030 34356 56082
rect 32396 55972 32452 55982
rect 32396 55878 32452 55916
rect 34300 55972 34356 56030
rect 31164 55298 31556 55300
rect 31164 55246 31166 55298
rect 31218 55246 31556 55298
rect 31164 55244 31556 55246
rect 31612 55524 31668 55534
rect 31164 54740 31220 55244
rect 30604 54226 30660 54236
rect 30828 54684 31220 54740
rect 30604 53732 30660 53742
rect 30828 53732 30884 54684
rect 30604 53730 30884 53732
rect 30604 53678 30606 53730
rect 30658 53678 30884 53730
rect 30604 53676 30884 53678
rect 30940 54514 30996 54526
rect 30940 54462 30942 54514
rect 30994 54462 30996 54514
rect 30604 53284 30660 53676
rect 30940 53508 30996 54462
rect 31500 54404 31556 54414
rect 31500 54310 31556 54348
rect 30940 53442 30996 53452
rect 31164 53844 31220 53854
rect 31164 53508 31220 53788
rect 31164 53442 31220 53452
rect 31612 53618 31668 55468
rect 31724 55412 31780 55422
rect 31780 55356 31892 55412
rect 31724 55346 31780 55356
rect 31724 55076 31780 55086
rect 31724 54982 31780 55020
rect 31836 54516 31892 55356
rect 32172 55300 32228 55310
rect 31724 54460 31892 54516
rect 32060 55298 32228 55300
rect 32060 55246 32174 55298
rect 32226 55246 32228 55298
rect 32060 55244 32228 55246
rect 31724 53732 31780 54460
rect 31836 54292 31892 54302
rect 31836 54198 31892 54236
rect 31724 53676 32004 53732
rect 31612 53566 31614 53618
rect 31666 53566 31668 53618
rect 31612 53396 31668 53566
rect 31724 53508 31780 53518
rect 31780 53452 31892 53508
rect 31724 53414 31780 53452
rect 31612 53330 31668 53340
rect 30604 53218 30660 53228
rect 31164 53172 31220 53182
rect 30716 53060 30772 53070
rect 30492 53004 30716 53060
rect 30380 52892 30548 52948
rect 29708 52108 29876 52164
rect 29484 51940 29540 51950
rect 29708 51940 29764 51950
rect 29372 51938 29652 51940
rect 29372 51886 29486 51938
rect 29538 51886 29652 51938
rect 29372 51884 29652 51886
rect 29484 51874 29540 51884
rect 29036 51716 29092 51726
rect 28700 51380 28756 51390
rect 28364 51378 28756 51380
rect 28364 51326 28702 51378
rect 28754 51326 28756 51378
rect 28364 51324 28756 51326
rect 28364 50818 28420 51324
rect 28700 51314 28756 51324
rect 29036 51378 29092 51660
rect 29036 51326 29038 51378
rect 29090 51326 29092 51378
rect 28364 50766 28366 50818
rect 28418 50766 28420 50818
rect 28364 50754 28420 50766
rect 29036 50428 29092 51326
rect 29372 51044 29428 51054
rect 29372 50708 29428 50988
rect 29484 50708 29540 50718
rect 29372 50706 29540 50708
rect 29372 50654 29486 50706
rect 29538 50654 29540 50706
rect 29372 50652 29540 50654
rect 29484 50642 29540 50652
rect 28252 49252 28308 49756
rect 28924 50372 29092 50428
rect 29372 50372 29428 50382
rect 28252 49186 28308 49196
rect 28364 49476 28420 49486
rect 28364 49028 28420 49420
rect 28924 49476 28980 50372
rect 28924 49410 28980 49420
rect 29260 50316 29372 50372
rect 28700 49084 29204 49140
rect 28364 48934 28420 48972
rect 28588 49028 28644 49038
rect 28476 48804 28532 48814
rect 28476 48710 28532 48748
rect 28252 48580 28308 48590
rect 28588 48580 28644 48972
rect 28700 49026 28756 49084
rect 28700 48974 28702 49026
rect 28754 48974 28756 49026
rect 28700 48962 28756 48974
rect 29148 49026 29204 49084
rect 29148 48974 29150 49026
rect 29202 48974 29204 49026
rect 29148 48962 29204 48974
rect 29260 49028 29316 50316
rect 29372 50306 29428 50316
rect 29596 50148 29652 51884
rect 29708 51846 29764 51884
rect 29820 51716 29876 52108
rect 30380 51940 30436 51950
rect 30380 51846 30436 51884
rect 29372 49812 29428 49822
rect 29596 49812 29652 50092
rect 29708 51660 29876 51716
rect 29708 50034 29764 51660
rect 29932 51604 29988 51614
rect 30156 51604 30212 51614
rect 29820 51492 29876 51502
rect 29932 51492 29988 51548
rect 29820 51490 29988 51492
rect 29820 51438 29822 51490
rect 29874 51438 29988 51490
rect 29820 51436 29988 51438
rect 30044 51548 30156 51604
rect 29820 51426 29876 51436
rect 30044 51268 30100 51548
rect 30156 51538 30212 51548
rect 29820 51212 30100 51268
rect 29820 51156 29876 51212
rect 29820 50818 29876 51100
rect 29820 50766 29822 50818
rect 29874 50766 29876 50818
rect 29820 50754 29876 50766
rect 30044 50932 30100 50942
rect 30044 50596 30100 50876
rect 30156 50820 30212 50830
rect 30156 50726 30212 50764
rect 30044 50482 30100 50540
rect 30044 50430 30046 50482
rect 30098 50430 30100 50482
rect 30044 50418 30100 50430
rect 30268 50596 30324 50606
rect 30268 50260 30324 50540
rect 29708 49982 29710 50034
rect 29762 49982 29764 50034
rect 29708 49970 29764 49982
rect 30044 50204 30324 50260
rect 29596 49756 29988 49812
rect 29372 49718 29428 49756
rect 29484 49700 29540 49710
rect 29484 49138 29540 49644
rect 29484 49086 29486 49138
rect 29538 49086 29540 49138
rect 29484 49074 29540 49086
rect 29372 49028 29428 49038
rect 29316 49026 29428 49028
rect 29316 48974 29374 49026
rect 29426 48974 29428 49026
rect 29316 48972 29428 48974
rect 29260 48934 29316 48972
rect 29372 48962 29428 48972
rect 29820 48914 29876 48926
rect 29820 48862 29822 48914
rect 29874 48862 29876 48914
rect 28252 47458 28308 48524
rect 28476 48524 28644 48580
rect 28812 48804 28868 48814
rect 28252 47406 28254 47458
rect 28306 47406 28308 47458
rect 28252 47124 28308 47406
rect 28364 48130 28420 48142
rect 28364 48078 28366 48130
rect 28418 48078 28420 48130
rect 28364 47460 28420 48078
rect 28476 47570 28532 48524
rect 28588 48132 28644 48142
rect 28588 48038 28644 48076
rect 28812 48020 28868 48748
rect 29036 48804 29092 48814
rect 28924 48020 28980 48030
rect 28812 48018 28980 48020
rect 28812 47966 28926 48018
rect 28978 47966 28980 48018
rect 28812 47964 28980 47966
rect 28476 47518 28478 47570
rect 28530 47518 28532 47570
rect 28476 47506 28532 47518
rect 28364 47394 28420 47404
rect 28252 47058 28308 47068
rect 28588 47346 28644 47358
rect 28588 47294 28590 47346
rect 28642 47294 28644 47346
rect 28364 46562 28420 46574
rect 28364 46510 28366 46562
rect 28418 46510 28420 46562
rect 27916 43538 28196 43540
rect 27916 43486 28030 43538
rect 28082 43486 28196 43538
rect 27916 43484 28196 43486
rect 28252 46004 28308 46014
rect 28252 43540 28308 45948
rect 28364 45220 28420 46510
rect 28588 46564 28644 47294
rect 28700 47012 28756 47022
rect 28756 46956 28868 47012
rect 28700 46946 28756 46956
rect 28588 46498 28644 46508
rect 28700 46676 28756 46686
rect 28588 46116 28644 46126
rect 28588 46002 28644 46060
rect 28588 45950 28590 46002
rect 28642 45950 28644 46002
rect 28588 45938 28644 45950
rect 28700 45780 28756 46620
rect 28700 45714 28756 45724
rect 28812 46676 28868 46956
rect 28924 46900 28980 47964
rect 28924 46834 28980 46844
rect 28924 46676 28980 46686
rect 28812 46674 28980 46676
rect 28812 46622 28926 46674
rect 28978 46622 28980 46674
rect 28812 46620 28980 46622
rect 28812 45556 28868 46620
rect 28924 46610 28980 46620
rect 28812 45490 28868 45500
rect 28924 45780 28980 45790
rect 28924 45330 28980 45724
rect 28924 45278 28926 45330
rect 28978 45278 28980 45330
rect 28924 45266 28980 45278
rect 28364 43764 28420 45164
rect 28476 45108 28532 45118
rect 28476 45014 28532 45052
rect 28700 45106 28756 45118
rect 28700 45054 28702 45106
rect 28754 45054 28756 45106
rect 28588 44548 28644 44558
rect 28588 44434 28644 44492
rect 28588 44382 28590 44434
rect 28642 44382 28644 44434
rect 28588 44370 28644 44382
rect 28700 44436 28756 45054
rect 28812 45108 28868 45118
rect 28812 45014 28868 45052
rect 29036 44772 29092 48748
rect 29596 48802 29652 48814
rect 29596 48750 29598 48802
rect 29650 48750 29652 48802
rect 29260 48692 29316 48702
rect 29260 48468 29316 48636
rect 29372 48468 29428 48478
rect 29260 48466 29428 48468
rect 29260 48414 29374 48466
rect 29426 48414 29428 48466
rect 29260 48412 29428 48414
rect 29372 48244 29428 48412
rect 29596 48468 29652 48750
rect 29820 48804 29876 48862
rect 29820 48738 29876 48748
rect 29596 48402 29652 48412
rect 29820 48468 29876 48478
rect 29820 48374 29876 48412
rect 29372 48178 29428 48188
rect 29596 47572 29652 47582
rect 29596 47478 29652 47516
rect 29148 47346 29204 47358
rect 29148 47294 29150 47346
rect 29202 47294 29204 47346
rect 29148 47124 29204 47294
rect 29148 47058 29204 47068
rect 29372 47346 29428 47358
rect 29372 47294 29374 47346
rect 29426 47294 29428 47346
rect 29260 46676 29316 46686
rect 29260 46582 29316 46620
rect 29260 46340 29316 46350
rect 29036 44706 29092 44716
rect 29148 45778 29204 45790
rect 29148 45726 29150 45778
rect 29202 45726 29204 45778
rect 29148 45106 29204 45726
rect 29260 45778 29316 46284
rect 29372 46004 29428 47294
rect 29708 47348 29764 47358
rect 29708 47254 29764 47292
rect 29820 47012 29876 47022
rect 29372 45938 29428 45948
rect 29484 46898 29540 46910
rect 29484 46846 29486 46898
rect 29538 46846 29540 46898
rect 29484 45892 29540 46846
rect 29596 46900 29652 46910
rect 29596 46786 29652 46844
rect 29596 46734 29598 46786
rect 29650 46734 29652 46786
rect 29596 46452 29652 46734
rect 29820 46786 29876 46956
rect 29820 46734 29822 46786
rect 29874 46734 29876 46786
rect 29820 46722 29876 46734
rect 29596 46386 29652 46396
rect 29932 46340 29988 49756
rect 30044 46900 30100 50204
rect 30380 49924 30436 49934
rect 30380 49830 30436 49868
rect 30156 49476 30212 49486
rect 30156 47124 30212 49420
rect 30268 48804 30324 48814
rect 30268 48710 30324 48748
rect 30492 48580 30548 52892
rect 30716 52946 30772 53004
rect 30716 52894 30718 52946
rect 30770 52894 30772 52946
rect 30716 52882 30772 52894
rect 30604 52162 30660 52174
rect 30604 52110 30606 52162
rect 30658 52110 30660 52162
rect 30604 51604 30660 52110
rect 30828 52164 30884 52174
rect 30828 52070 30884 52108
rect 31164 52162 31220 53116
rect 31836 52724 31892 53452
rect 31948 53172 32004 53676
rect 31948 53078 32004 53116
rect 31836 52658 31892 52668
rect 32060 52612 32116 55244
rect 32172 55234 32228 55244
rect 33852 55298 33908 55310
rect 33852 55246 33854 55298
rect 33906 55246 33908 55298
rect 32732 55188 32788 55198
rect 33068 55188 33124 55198
rect 32732 55094 32788 55132
rect 32956 55186 33124 55188
rect 32956 55134 33070 55186
rect 33122 55134 33124 55186
rect 32956 55132 33124 55134
rect 32284 53730 32340 53742
rect 32284 53678 32286 53730
rect 32338 53678 32340 53730
rect 32172 53620 32228 53630
rect 32172 53526 32228 53564
rect 32284 53396 32340 53678
rect 32956 53732 33012 55132
rect 33068 55122 33124 55132
rect 33180 55188 33236 55198
rect 33180 55076 33236 55132
rect 33404 55076 33460 55086
rect 33180 55074 33348 55076
rect 33180 55022 33182 55074
rect 33234 55022 33348 55074
rect 33180 55020 33348 55022
rect 33180 55010 33236 55020
rect 33180 53956 33236 53966
rect 32956 53666 33012 53676
rect 33068 53730 33124 53742
rect 33068 53678 33070 53730
rect 33122 53678 33124 53730
rect 32060 52546 32116 52556
rect 32172 53340 32340 53396
rect 32172 52388 32228 53340
rect 33068 53284 33124 53678
rect 33180 53506 33236 53900
rect 33292 53620 33348 55020
rect 33404 55074 33572 55076
rect 33404 55022 33406 55074
rect 33458 55022 33572 55074
rect 33404 55020 33572 55022
rect 33404 55010 33460 55020
rect 33292 53554 33348 53564
rect 33180 53454 33182 53506
rect 33234 53454 33236 53506
rect 33180 53442 33236 53454
rect 33068 53228 33460 53284
rect 32284 53172 32340 53182
rect 33068 53172 33124 53228
rect 32284 53170 33124 53172
rect 32284 53118 32286 53170
rect 32338 53118 33124 53170
rect 32284 53116 33124 53118
rect 32284 53106 32340 53116
rect 33180 52836 33236 52846
rect 33068 52834 33236 52836
rect 33068 52782 33182 52834
rect 33234 52782 33236 52834
rect 33068 52780 33236 52782
rect 32956 52724 33012 52734
rect 32732 52722 33012 52724
rect 32732 52670 32958 52722
rect 33010 52670 33012 52722
rect 32732 52668 33012 52670
rect 32172 52332 32340 52388
rect 31836 52276 31892 52286
rect 31836 52182 31892 52220
rect 31164 52110 31166 52162
rect 31218 52110 31220 52162
rect 31164 52098 31220 52110
rect 32172 52162 32228 52174
rect 32172 52110 32174 52162
rect 32226 52110 32228 52162
rect 30604 51538 30660 51548
rect 31164 51604 31220 51614
rect 31724 51604 31780 51614
rect 31164 51602 31780 51604
rect 31164 51550 31166 51602
rect 31218 51550 31726 51602
rect 31778 51550 31780 51602
rect 31164 51548 31780 51550
rect 31164 51538 31220 51548
rect 31724 51538 31780 51548
rect 30716 51378 30772 51390
rect 30716 51326 30718 51378
rect 30770 51326 30772 51378
rect 30716 50820 30772 51326
rect 30716 50754 30772 50764
rect 30940 51378 30996 51390
rect 30940 51326 30942 51378
rect 30994 51326 30996 51378
rect 30940 50706 30996 51326
rect 31276 51380 31332 51390
rect 32172 51380 32228 52110
rect 32284 51492 32340 52332
rect 32732 52162 32788 52668
rect 32956 52658 33012 52668
rect 33068 52724 33124 52780
rect 33180 52770 33236 52780
rect 32732 52110 32734 52162
rect 32786 52110 32788 52162
rect 32284 51436 32452 51492
rect 31276 51286 31332 51324
rect 31724 51324 32228 51380
rect 31164 51266 31220 51278
rect 31164 51214 31166 51266
rect 31218 51214 31220 51266
rect 31164 50820 31220 51214
rect 31164 50754 31220 50764
rect 31612 51044 31668 51054
rect 30940 50654 30942 50706
rect 30994 50654 30996 50706
rect 30940 50642 30996 50654
rect 30828 50596 30884 50606
rect 30716 50594 30884 50596
rect 30716 50542 30830 50594
rect 30882 50542 30884 50594
rect 30716 50540 30884 50542
rect 30604 50484 30660 50494
rect 30604 50370 30660 50428
rect 30716 50428 30772 50540
rect 30828 50530 30884 50540
rect 31052 50596 31108 50606
rect 31052 50502 31108 50540
rect 31388 50484 31444 50522
rect 30716 50372 30884 50428
rect 31388 50418 31444 50428
rect 31612 50482 31668 50988
rect 31724 50818 31780 51324
rect 32284 51266 32340 51278
rect 32284 51214 32286 51266
rect 32338 51214 32340 51266
rect 32060 51156 32116 51166
rect 32060 51062 32116 51100
rect 32284 51044 32340 51214
rect 32284 50978 32340 50988
rect 31724 50766 31726 50818
rect 31778 50766 31780 50818
rect 31724 50754 31780 50766
rect 32284 50708 32340 50718
rect 32284 50594 32340 50652
rect 32284 50542 32286 50594
rect 32338 50542 32340 50594
rect 32284 50530 32340 50542
rect 31612 50430 31614 50482
rect 31666 50430 31668 50482
rect 31612 50418 31668 50430
rect 32172 50484 32228 50494
rect 32396 50484 32452 51436
rect 32732 50484 32788 52110
rect 32956 51604 33012 51614
rect 32956 50818 33012 51548
rect 32956 50766 32958 50818
rect 33010 50766 33012 50818
rect 32956 50754 33012 50766
rect 32396 50428 32564 50484
rect 30604 50318 30606 50370
rect 30658 50318 30660 50370
rect 30604 48804 30660 50318
rect 30716 50260 30772 50270
rect 30716 49138 30772 50204
rect 30716 49086 30718 49138
rect 30770 49086 30772 49138
rect 30716 49028 30772 49086
rect 30828 49812 30884 50372
rect 31724 50148 31780 50158
rect 31612 50092 31724 50148
rect 31612 50034 31668 50092
rect 31724 50082 31780 50092
rect 31612 49982 31614 50034
rect 31666 49982 31668 50034
rect 31612 49970 31668 49982
rect 31276 49924 31332 49934
rect 31500 49924 31556 49934
rect 31276 49830 31332 49868
rect 31388 49922 31556 49924
rect 31388 49870 31502 49922
rect 31554 49870 31556 49922
rect 31388 49868 31556 49870
rect 30828 49140 30884 49756
rect 31388 49812 31444 49868
rect 31500 49858 31556 49868
rect 31388 49746 31444 49756
rect 31724 49810 31780 49822
rect 31724 49758 31726 49810
rect 31778 49758 31780 49810
rect 31724 49588 31780 49758
rect 31052 49532 31780 49588
rect 31836 49810 31892 49822
rect 31836 49758 31838 49810
rect 31890 49758 31892 49810
rect 30828 49074 30884 49084
rect 30940 49476 30996 49486
rect 30716 48962 30772 48972
rect 30604 48748 30884 48804
rect 30492 48524 30772 48580
rect 30268 48468 30324 48478
rect 30324 48412 30436 48468
rect 30268 48402 30324 48412
rect 30268 48244 30324 48254
rect 30268 48150 30324 48188
rect 30380 48020 30436 48412
rect 30156 47058 30212 47068
rect 30268 47964 30436 48020
rect 30604 48354 30660 48366
rect 30604 48302 30606 48354
rect 30658 48302 30660 48354
rect 30044 46834 30100 46844
rect 30156 46788 30212 46798
rect 30156 46694 30212 46732
rect 30268 46674 30324 47964
rect 30492 47684 30548 47694
rect 30492 47590 30548 47628
rect 30380 47348 30436 47358
rect 30604 47348 30660 48302
rect 30436 47292 30660 47348
rect 30380 47254 30436 47292
rect 30268 46622 30270 46674
rect 30322 46622 30324 46674
rect 30268 46610 30324 46622
rect 29932 46274 29988 46284
rect 30268 46340 30324 46350
rect 30044 46004 30100 46014
rect 30044 45910 30100 45948
rect 29484 45826 29540 45836
rect 30156 45890 30212 45902
rect 30156 45838 30158 45890
rect 30210 45838 30212 45890
rect 29260 45726 29262 45778
rect 29314 45726 29316 45778
rect 29260 45714 29316 45726
rect 29484 45668 29540 45678
rect 29484 45666 30100 45668
rect 29484 45614 29486 45666
rect 29538 45614 30100 45666
rect 29484 45612 30100 45614
rect 29484 45602 29540 45612
rect 29260 45556 29316 45566
rect 29316 45500 29428 45556
rect 29260 45490 29316 45500
rect 29372 45220 29428 45500
rect 29932 45444 29988 45454
rect 29484 45220 29540 45230
rect 29372 45218 29540 45220
rect 29372 45166 29486 45218
rect 29538 45166 29540 45218
rect 29372 45164 29540 45166
rect 29484 45154 29540 45164
rect 29708 45220 29764 45230
rect 29708 45126 29764 45164
rect 29148 45054 29150 45106
rect 29202 45054 29204 45106
rect 28700 44370 28756 44380
rect 29148 43876 29204 45054
rect 29596 44994 29652 45006
rect 29596 44942 29598 44994
rect 29650 44942 29652 44994
rect 29596 44772 29652 44942
rect 29372 44716 29652 44772
rect 29260 44548 29316 44558
rect 29260 44454 29316 44492
rect 29372 44436 29428 44716
rect 29372 44370 29428 44380
rect 29484 44324 29540 44334
rect 29148 43820 29316 43876
rect 28364 43708 28532 43764
rect 28252 43484 28420 43540
rect 27580 42662 27636 42700
rect 27692 43428 27748 43438
rect 27916 43428 27972 43484
rect 28028 43474 28084 43484
rect 27692 43426 27972 43428
rect 27692 43374 27694 43426
rect 27746 43374 27972 43426
rect 27692 43372 27972 43374
rect 27356 42140 27524 42196
rect 26460 41570 26516 41580
rect 26348 41188 26404 41356
rect 26236 41132 26404 41188
rect 26236 41074 26292 41132
rect 26684 41076 26740 41086
rect 26236 41022 26238 41074
rect 26290 41022 26292 41074
rect 26236 41010 26292 41022
rect 26348 41074 26740 41076
rect 26348 41022 26686 41074
rect 26738 41022 26740 41074
rect 26348 41020 26740 41022
rect 26124 40964 26180 40974
rect 26124 40870 26180 40908
rect 25676 40684 25844 40740
rect 25676 40402 25732 40684
rect 25676 40350 25678 40402
rect 25730 40350 25732 40402
rect 25452 39554 25508 39564
rect 25564 40292 25620 40302
rect 25340 39442 25396 39452
rect 25228 38612 25508 38668
rect 24948 38556 25172 38612
rect 24892 38546 24948 38556
rect 24556 38162 24836 38164
rect 24556 38110 24558 38162
rect 24610 38110 24836 38162
rect 24556 38108 24836 38110
rect 24556 38098 24612 38108
rect 24780 38050 24836 38108
rect 24780 37998 24782 38050
rect 24834 37998 24836 38050
rect 24780 37986 24836 37998
rect 25116 38052 25172 38556
rect 25228 38052 25284 38062
rect 25116 38050 25284 38052
rect 25116 37998 25230 38050
rect 25282 37998 25284 38050
rect 25116 37996 25284 37998
rect 25228 37986 25284 37996
rect 25452 38050 25508 38612
rect 25452 37998 25454 38050
rect 25506 37998 25508 38050
rect 25452 37986 25508 37998
rect 23996 37938 24164 37940
rect 23996 37886 23998 37938
rect 24050 37886 24164 37938
rect 23996 37884 24164 37886
rect 23996 37874 24052 37884
rect 24220 37828 24276 37838
rect 23996 37492 24052 37502
rect 23996 37398 24052 37436
rect 24220 37378 24276 37772
rect 25340 37826 25396 37838
rect 25340 37774 25342 37826
rect 25394 37774 25396 37826
rect 24332 37492 24388 37502
rect 24332 37398 24388 37436
rect 24220 37326 24222 37378
rect 24274 37326 24276 37378
rect 24220 37314 24276 37326
rect 25340 37380 25396 37774
rect 25340 37314 25396 37324
rect 24556 37268 24612 37278
rect 24556 37266 24724 37268
rect 24556 37214 24558 37266
rect 24610 37214 24724 37266
rect 24556 37212 24724 37214
rect 24556 37202 24612 37212
rect 24668 36596 24724 37212
rect 24668 36540 25284 36596
rect 23996 36482 24052 36494
rect 23996 36430 23998 36482
rect 24050 36430 24052 36482
rect 23996 36372 24052 36430
rect 24668 36482 24724 36540
rect 24668 36430 24670 36482
rect 24722 36430 24724 36482
rect 24668 36418 24724 36430
rect 23996 36306 24052 36316
rect 24332 36370 24388 36382
rect 24332 36318 24334 36370
rect 24386 36318 24388 36370
rect 23884 36092 24276 36148
rect 23716 34300 23828 34356
rect 24220 34914 24276 36092
rect 24332 35924 24388 36318
rect 24892 36370 24948 36382
rect 24892 36318 24894 36370
rect 24946 36318 24948 36370
rect 24332 35858 24388 35868
rect 24668 36036 24724 36046
rect 24668 35922 24724 35980
rect 24668 35870 24670 35922
rect 24722 35870 24724 35922
rect 24668 35858 24724 35870
rect 24220 34862 24222 34914
rect 24274 34862 24276 34914
rect 23660 34290 23716 34300
rect 24220 34020 24276 34862
rect 24220 33954 24276 33964
rect 24780 34916 24836 34926
rect 23436 33460 23492 33516
rect 24668 33572 24724 33582
rect 24780 33572 24836 34860
rect 24892 34468 24948 36318
rect 25228 35810 25284 36540
rect 25564 36482 25620 40236
rect 25676 39060 25732 40350
rect 25788 40404 25844 40414
rect 25788 40310 25844 40348
rect 26012 39844 26068 39854
rect 26012 39730 26068 39788
rect 26012 39678 26014 39730
rect 26066 39678 26068 39730
rect 26012 39666 26068 39678
rect 25676 38994 25732 39004
rect 26012 39060 26068 39070
rect 26012 38052 26068 39004
rect 25564 36430 25566 36482
rect 25618 36430 25620 36482
rect 25340 36036 25396 36046
rect 25340 35922 25396 35980
rect 25340 35870 25342 35922
rect 25394 35870 25396 35922
rect 25340 35858 25396 35870
rect 25564 35924 25620 36430
rect 25900 37996 26068 38052
rect 26124 38836 26180 38846
rect 25676 36260 25732 36270
rect 25676 36166 25732 36204
rect 25564 35868 25732 35924
rect 25228 35758 25230 35810
rect 25282 35758 25284 35810
rect 25228 35746 25284 35758
rect 25564 35698 25620 35710
rect 25564 35646 25566 35698
rect 25618 35646 25620 35698
rect 25564 34804 25620 35646
rect 25676 35474 25732 35868
rect 25676 35422 25678 35474
rect 25730 35422 25732 35474
rect 25676 35410 25732 35422
rect 25900 35028 25956 37996
rect 26012 37828 26068 37838
rect 26012 37734 26068 37772
rect 26012 35586 26068 35598
rect 26012 35534 26014 35586
rect 26066 35534 26068 35586
rect 26012 35474 26068 35534
rect 26012 35422 26014 35474
rect 26066 35422 26068 35474
rect 26012 35410 26068 35422
rect 26124 35364 26180 38780
rect 26236 38276 26292 38286
rect 26236 38050 26292 38220
rect 26236 37998 26238 38050
rect 26290 37998 26292 38050
rect 26236 37604 26292 37998
rect 26236 37538 26292 37548
rect 26236 36708 26292 36718
rect 26348 36708 26404 41020
rect 26684 41010 26740 41020
rect 26796 40964 26852 42140
rect 27468 42084 27524 42140
rect 27468 42082 27636 42084
rect 27468 42030 27470 42082
rect 27522 42030 27636 42082
rect 27468 42028 27636 42030
rect 27468 42018 27524 42028
rect 27356 41972 27412 41982
rect 27356 41878 27412 41916
rect 27020 41860 27076 41870
rect 27020 41186 27076 41804
rect 27020 41134 27022 41186
rect 27074 41134 27076 41186
rect 27020 41122 27076 41134
rect 27356 40964 27412 40974
rect 26796 40962 27412 40964
rect 26796 40910 26798 40962
rect 26850 40910 27358 40962
rect 27410 40910 27412 40962
rect 26796 40908 27412 40910
rect 26572 40628 26628 40638
rect 26572 40534 26628 40572
rect 26796 39060 26852 40908
rect 27356 40898 27412 40908
rect 27132 40516 27188 40526
rect 27356 40516 27412 40526
rect 27188 40514 27412 40516
rect 27188 40462 27358 40514
rect 27410 40462 27412 40514
rect 27188 40460 27412 40462
rect 27132 40422 27188 40460
rect 27356 40450 27412 40460
rect 27244 40292 27300 40302
rect 26796 38994 26852 39004
rect 26908 39396 26964 39406
rect 26572 38052 26628 38062
rect 26908 38052 26964 39340
rect 27244 38668 27300 40236
rect 27580 39844 27636 42028
rect 27692 41076 27748 43372
rect 28252 43314 28308 43326
rect 28252 43262 28254 43314
rect 28306 43262 28308 43314
rect 27804 43092 27860 43102
rect 27804 41972 27860 43036
rect 28028 42978 28084 42990
rect 28028 42926 28030 42978
rect 28082 42926 28084 42978
rect 27916 42420 27972 42430
rect 27916 42194 27972 42364
rect 27916 42142 27918 42194
rect 27970 42142 27972 42194
rect 27916 42130 27972 42142
rect 27804 41916 27972 41972
rect 27804 41412 27860 41422
rect 27804 41298 27860 41356
rect 27804 41246 27806 41298
rect 27858 41246 27860 41298
rect 27804 41234 27860 41246
rect 27692 41020 27860 41076
rect 27692 40514 27748 40526
rect 27692 40462 27694 40514
rect 27746 40462 27748 40514
rect 27692 40292 27748 40462
rect 27692 40226 27748 40236
rect 27580 39778 27636 39788
rect 27692 39732 27748 39742
rect 27692 39618 27748 39676
rect 27692 39566 27694 39618
rect 27746 39566 27748 39618
rect 27692 39554 27748 39566
rect 27132 38612 27300 38668
rect 27468 38836 27524 38846
rect 27132 38276 27188 38612
rect 26572 37958 26628 37996
rect 26684 37996 26964 38052
rect 27020 38220 27188 38276
rect 26572 37604 26628 37614
rect 26572 36932 26628 37548
rect 26684 37044 26740 37996
rect 26796 37826 26852 37838
rect 26796 37774 26798 37826
rect 26850 37774 26852 37826
rect 26796 37716 26852 37774
rect 26908 37828 26964 37838
rect 26908 37734 26964 37772
rect 26796 37650 26852 37660
rect 26908 37380 26964 37390
rect 26908 37266 26964 37324
rect 26908 37214 26910 37266
rect 26962 37214 26964 37266
rect 26908 37202 26964 37214
rect 27020 37156 27076 38220
rect 27132 38050 27188 38062
rect 27132 37998 27134 38050
rect 27186 37998 27188 38050
rect 27132 37940 27188 37998
rect 27132 37874 27188 37884
rect 27356 37826 27412 37838
rect 27356 37774 27358 37826
rect 27410 37774 27412 37826
rect 27244 37266 27300 37278
rect 27244 37214 27246 37266
rect 27298 37214 27300 37266
rect 27020 37100 27188 37156
rect 26684 36988 27076 37044
rect 26572 36876 26852 36932
rect 26292 36652 26404 36708
rect 26236 36614 26292 36652
rect 26572 36596 26628 36606
rect 26572 36502 26628 36540
rect 26460 36484 26516 36494
rect 26460 36370 26516 36428
rect 26460 36318 26462 36370
rect 26514 36318 26516 36370
rect 26460 36306 26516 36318
rect 26684 36260 26740 36270
rect 26684 36036 26740 36204
rect 26796 36148 26852 36876
rect 27020 36258 27076 36988
rect 27132 36708 27188 37100
rect 27244 36820 27300 37214
rect 27356 37268 27412 37774
rect 27468 37490 27524 38780
rect 27804 38834 27860 41020
rect 27916 40628 27972 41916
rect 27916 40562 27972 40572
rect 28028 40404 28084 42926
rect 28252 42532 28308 43262
rect 28252 42466 28308 42476
rect 28140 42082 28196 42094
rect 28140 42030 28142 42082
rect 28194 42030 28196 42082
rect 28140 40628 28196 42030
rect 28364 41972 28420 43484
rect 28476 43092 28532 43708
rect 28700 43708 29092 43764
rect 28588 43652 28644 43662
rect 28700 43652 28756 43708
rect 28644 43596 28756 43652
rect 29036 43650 29092 43708
rect 29036 43598 29038 43650
rect 29090 43598 29092 43650
rect 28588 43586 28644 43596
rect 29036 43586 29092 43598
rect 29148 43652 29204 43662
rect 29148 43558 29204 43596
rect 29260 43428 29316 43820
rect 29148 43372 29316 43428
rect 28588 43316 28644 43326
rect 28588 43222 28644 43260
rect 29036 43314 29092 43326
rect 29036 43262 29038 43314
rect 29090 43262 29092 43314
rect 28924 43204 28980 43214
rect 28476 43036 28644 43092
rect 28364 41906 28420 41916
rect 28476 41972 28532 41982
rect 28588 41972 28644 43036
rect 28700 42756 28756 42766
rect 28924 42756 28980 43148
rect 29036 43092 29092 43262
rect 29036 43026 29092 43036
rect 29036 42756 29092 42766
rect 28924 42754 29092 42756
rect 28924 42702 29038 42754
rect 29090 42702 29092 42754
rect 28924 42700 29092 42702
rect 28700 42662 28756 42700
rect 29036 42690 29092 42700
rect 28924 42084 28980 42094
rect 28924 41990 28980 42028
rect 29148 42082 29204 43372
rect 29372 42644 29428 42654
rect 29148 42030 29150 42082
rect 29202 42030 29204 42082
rect 28476 41970 28644 41972
rect 28476 41918 28478 41970
rect 28530 41918 28644 41970
rect 28476 41916 28644 41918
rect 28476 41906 28532 41916
rect 28476 41748 28532 41758
rect 28364 40628 28420 40638
rect 28140 40572 28308 40628
rect 27916 40402 28084 40404
rect 27916 40350 28030 40402
rect 28082 40350 28084 40402
rect 27916 40348 28084 40350
rect 27916 39618 27972 40348
rect 28028 40338 28084 40348
rect 27916 39566 27918 39618
rect 27970 39566 27972 39618
rect 27916 39554 27972 39566
rect 28028 39732 28084 39742
rect 28028 39396 28084 39676
rect 28028 39330 28084 39340
rect 27804 38782 27806 38834
rect 27858 38782 27860 38834
rect 27804 38668 27860 38782
rect 28252 38668 28308 40572
rect 28364 40514 28420 40572
rect 28364 40462 28366 40514
rect 28418 40462 28420 40514
rect 28364 40450 28420 40462
rect 28476 38946 28532 41692
rect 28588 40516 28644 41916
rect 28700 41076 28756 41086
rect 28700 40982 28756 41020
rect 29036 40964 29092 40974
rect 28588 40422 28644 40460
rect 28700 40626 28756 40638
rect 28700 40574 28702 40626
rect 28754 40574 28756 40626
rect 28588 39396 28644 39406
rect 28588 39302 28644 39340
rect 28476 38894 28478 38946
rect 28530 38894 28532 38946
rect 28476 38882 28532 38894
rect 28700 38668 28756 40574
rect 27692 38610 27748 38622
rect 27804 38612 28196 38668
rect 28252 38612 28420 38668
rect 27692 38558 27694 38610
rect 27746 38558 27748 38610
rect 27692 37940 27748 38558
rect 27916 38162 27972 38174
rect 27916 38110 27918 38162
rect 27970 38110 27972 38162
rect 27692 37884 27860 37940
rect 27468 37438 27470 37490
rect 27522 37438 27524 37490
rect 27468 37426 27524 37438
rect 27692 37716 27748 37726
rect 27580 37268 27636 37278
rect 27692 37268 27748 37660
rect 27804 37492 27860 37884
rect 27804 37426 27860 37436
rect 27356 37212 27524 37268
rect 27468 37044 27524 37212
rect 27580 37266 27748 37268
rect 27580 37214 27582 37266
rect 27634 37214 27748 37266
rect 27580 37212 27748 37214
rect 27804 37266 27860 37278
rect 27804 37214 27806 37266
rect 27858 37214 27860 37266
rect 27580 37202 27636 37212
rect 27468 36978 27524 36988
rect 27804 37044 27860 37214
rect 27804 36978 27860 36988
rect 27916 36932 27972 38110
rect 28140 38164 28196 38612
rect 28140 37938 28196 38108
rect 28140 37886 28142 37938
rect 28194 37886 28196 37938
rect 28140 37874 28196 37886
rect 28252 37940 28308 37950
rect 28028 37828 28084 37838
rect 28028 37716 28084 37772
rect 28028 37660 28196 37716
rect 28140 37266 28196 37660
rect 28252 37490 28308 37884
rect 28252 37438 28254 37490
rect 28306 37438 28308 37490
rect 28252 37426 28308 37438
rect 28140 37214 28142 37266
rect 28194 37214 28196 37266
rect 28140 37202 28196 37214
rect 27916 36876 28084 36932
rect 27244 36764 27636 36820
rect 27580 36708 27636 36764
rect 27132 36652 27524 36708
rect 27580 36652 27972 36708
rect 27356 36482 27412 36494
rect 27356 36430 27358 36482
rect 27410 36430 27412 36482
rect 27356 36372 27412 36430
rect 27356 36306 27412 36316
rect 27020 36206 27022 36258
rect 27074 36206 27076 36258
rect 27020 36194 27076 36206
rect 26796 36092 26964 36148
rect 26684 35970 26740 35980
rect 26908 35810 26964 36092
rect 27356 36036 27412 36046
rect 27020 35924 27076 35934
rect 27244 35924 27300 35934
rect 27356 35924 27412 35980
rect 27020 35922 27188 35924
rect 27020 35870 27022 35922
rect 27074 35870 27188 35922
rect 27020 35868 27188 35870
rect 27020 35858 27076 35868
rect 26908 35758 26910 35810
rect 26962 35758 26964 35810
rect 26908 35746 26964 35758
rect 27132 35700 27188 35868
rect 27244 35922 27412 35924
rect 27244 35870 27246 35922
rect 27298 35870 27412 35922
rect 27244 35868 27412 35870
rect 27244 35858 27300 35868
rect 27356 35700 27412 35710
rect 27132 35644 27356 35700
rect 26348 35364 26404 35374
rect 26124 35308 26348 35364
rect 26348 35298 26404 35308
rect 25900 34934 25956 34972
rect 26684 35028 26740 35038
rect 26348 34916 26404 34926
rect 26348 34822 26404 34860
rect 25564 34738 25620 34748
rect 26684 34802 26740 34972
rect 27356 35026 27412 35644
rect 27356 34974 27358 35026
rect 27410 34974 27412 35026
rect 27356 34962 27412 34974
rect 26684 34750 26686 34802
rect 26738 34750 26740 34802
rect 26684 34738 26740 34750
rect 27244 34916 27300 34926
rect 27244 34804 27300 34860
rect 27468 34804 27524 36652
rect 27580 36484 27636 36494
rect 27580 36390 27636 36428
rect 27916 36482 27972 36652
rect 27916 36430 27918 36482
rect 27970 36430 27972 36482
rect 27916 36418 27972 36430
rect 27244 34748 27636 34804
rect 24892 34402 24948 34412
rect 26012 34356 26068 34366
rect 25788 34354 26068 34356
rect 25788 34302 26014 34354
rect 26066 34302 26068 34354
rect 25788 34300 26068 34302
rect 25676 34244 25732 34254
rect 25564 34132 25620 34142
rect 25564 34038 25620 34076
rect 25676 33908 25732 34188
rect 25676 33842 25732 33852
rect 25788 33684 25844 34300
rect 26012 34290 26068 34300
rect 26236 34356 26292 34366
rect 26236 34262 26292 34300
rect 25900 34132 25956 34142
rect 26348 34132 26404 34142
rect 25900 34130 26180 34132
rect 25900 34078 25902 34130
rect 25954 34078 26180 34130
rect 25900 34076 26180 34078
rect 25900 34066 25956 34076
rect 25228 33628 25844 33684
rect 26012 33908 26068 33918
rect 24668 33570 24836 33572
rect 24668 33518 24670 33570
rect 24722 33518 24836 33570
rect 24668 33516 24836 33518
rect 25004 33572 25060 33582
rect 24668 33506 24724 33516
rect 23548 33460 23604 33470
rect 23436 33458 23604 33460
rect 23436 33406 23550 33458
rect 23602 33406 23604 33458
rect 23436 33404 23604 33406
rect 21980 33348 22036 33358
rect 21980 33254 22036 33292
rect 22652 33348 22708 33358
rect 22652 33346 22820 33348
rect 22652 33294 22654 33346
rect 22706 33294 22820 33346
rect 22652 33292 22820 33294
rect 22652 33282 22708 33292
rect 22092 33236 22148 33246
rect 22092 33142 22148 33180
rect 22204 33122 22260 33134
rect 22204 33070 22206 33122
rect 22258 33070 22260 33122
rect 22204 32564 22260 33070
rect 22764 32786 22820 33292
rect 22988 32788 23044 33404
rect 23548 33394 23604 33404
rect 24332 33460 24388 33470
rect 23996 33124 24052 33134
rect 23996 33030 24052 33068
rect 24332 33122 24388 33404
rect 24444 33346 24500 33358
rect 24444 33294 24446 33346
rect 24498 33294 24500 33346
rect 24444 33236 24500 33294
rect 25004 33346 25060 33516
rect 25228 33570 25284 33628
rect 25228 33518 25230 33570
rect 25282 33518 25284 33570
rect 25228 33506 25284 33518
rect 25004 33294 25006 33346
rect 25058 33294 25060 33346
rect 25004 33282 25060 33294
rect 25676 33348 25732 33358
rect 25676 33254 25732 33292
rect 25900 33346 25956 33358
rect 25900 33294 25902 33346
rect 25954 33294 25956 33346
rect 24444 33170 24500 33180
rect 25564 33236 25620 33246
rect 24332 33070 24334 33122
rect 24386 33070 24388 33122
rect 24332 33058 24388 33070
rect 24780 33124 24836 33134
rect 22764 32734 22766 32786
rect 22818 32734 22820 32786
rect 22764 32722 22820 32734
rect 22876 32786 23044 32788
rect 22876 32734 22990 32786
rect 23042 32734 23044 32786
rect 22876 32732 23044 32734
rect 22652 32564 22708 32574
rect 22876 32564 22932 32732
rect 22988 32722 23044 32732
rect 24780 32786 24836 33068
rect 24780 32734 24782 32786
rect 24834 32734 24836 32786
rect 24780 32722 24836 32734
rect 25452 33124 25508 33134
rect 25452 32786 25508 33068
rect 25452 32734 25454 32786
rect 25506 32734 25508 32786
rect 25452 32722 25508 32734
rect 23436 32676 23492 32686
rect 23436 32582 23492 32620
rect 25228 32676 25284 32686
rect 25228 32582 25284 32620
rect 22204 32562 22932 32564
rect 22204 32510 22654 32562
rect 22706 32510 22932 32562
rect 22204 32508 22932 32510
rect 23100 32562 23156 32574
rect 23100 32510 23102 32562
rect 23154 32510 23156 32562
rect 22652 32498 22708 32508
rect 23100 32340 23156 32510
rect 25564 32450 25620 33180
rect 25900 33124 25956 33294
rect 26012 33348 26068 33852
rect 26124 33684 26180 34076
rect 26348 33908 26404 34076
rect 26348 33852 26628 33908
rect 26236 33740 26516 33796
rect 26236 33684 26292 33740
rect 26124 33628 26292 33684
rect 26348 33570 26404 33582
rect 26348 33518 26350 33570
rect 26402 33518 26404 33570
rect 26236 33348 26292 33358
rect 26012 33346 26292 33348
rect 26012 33294 26238 33346
rect 26290 33294 26292 33346
rect 26012 33292 26292 33294
rect 26236 33282 26292 33292
rect 25900 33058 25956 33068
rect 25788 32564 25844 32574
rect 25788 32562 25956 32564
rect 25788 32510 25790 32562
rect 25842 32510 25956 32562
rect 25788 32508 25956 32510
rect 25788 32498 25844 32508
rect 25564 32398 25566 32450
rect 25618 32398 25620 32450
rect 25564 32386 25620 32398
rect 23100 32274 23156 32284
rect 23548 32340 23604 32350
rect 23548 32246 23604 32284
rect 24220 32340 24276 32350
rect 21196 31826 21252 31836
rect 21980 31780 22036 31790
rect 21308 31666 21364 31678
rect 21308 31614 21310 31666
rect 21362 31614 21364 31666
rect 21308 30772 21364 31614
rect 21980 31554 22036 31724
rect 21980 31502 21982 31554
rect 22034 31502 22036 31554
rect 21980 31490 22036 31502
rect 21868 31108 21924 31118
rect 21868 31014 21924 31052
rect 21308 30706 21364 30716
rect 21756 30884 21812 30894
rect 21756 30322 21812 30828
rect 23996 30772 24052 30782
rect 24052 30716 24164 30772
rect 23996 30706 24052 30716
rect 21756 30270 21758 30322
rect 21810 30270 21812 30322
rect 21756 30258 21812 30270
rect 23996 30322 24052 30334
rect 23996 30270 23998 30322
rect 24050 30270 24052 30322
rect 21980 30212 22036 30222
rect 22316 30212 22372 30222
rect 21980 30210 22148 30212
rect 21980 30158 21982 30210
rect 22034 30158 22148 30210
rect 21980 30156 22148 30158
rect 21980 30146 22036 30156
rect 21308 30100 21364 30110
rect 21308 30006 21364 30044
rect 21532 29988 21588 29998
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20636 29810 20692 29820
rect 21420 29986 21588 29988
rect 21420 29934 21534 29986
rect 21586 29934 21588 29986
rect 21420 29932 21588 29934
rect 19836 29754 20100 29764
rect 19964 29652 20020 29662
rect 19964 29558 20020 29596
rect 20636 29652 20692 29662
rect 19852 29540 19908 29550
rect 19628 29484 19852 29540
rect 19852 29446 19908 29484
rect 18844 29428 18900 29438
rect 18732 29426 18900 29428
rect 18732 29374 18846 29426
rect 18898 29374 18900 29426
rect 18732 29372 18900 29374
rect 17724 29148 18228 29204
rect 17612 28578 17668 28588
rect 17836 28642 17892 28654
rect 17836 28590 17838 28642
rect 17890 28590 17892 28642
rect 17612 28420 17668 28430
rect 17836 28420 17892 28590
rect 18172 28530 18228 29148
rect 18508 29138 18564 29148
rect 18620 29314 18676 29326
rect 18620 29262 18622 29314
rect 18674 29262 18676 29314
rect 18620 28980 18676 29262
rect 18620 28914 18676 28924
rect 18620 28756 18676 28766
rect 18732 28756 18788 29372
rect 18844 29362 18900 29372
rect 18956 29316 19012 29326
rect 18956 29222 19012 29260
rect 19740 29316 19796 29326
rect 19740 29222 19796 29260
rect 18172 28478 18174 28530
rect 18226 28478 18228 28530
rect 18172 28466 18228 28478
rect 18396 28754 18788 28756
rect 18396 28702 18622 28754
rect 18674 28702 18788 28754
rect 18396 28700 18788 28702
rect 19292 28868 19348 28878
rect 19292 28754 19348 28812
rect 19292 28702 19294 28754
rect 19346 28702 19348 28754
rect 17612 28418 17892 28420
rect 17612 28366 17614 28418
rect 17666 28366 17892 28418
rect 17612 28364 17892 28366
rect 17612 27972 17668 28364
rect 17612 27906 17668 27916
rect 17388 27860 17444 27870
rect 17388 27766 17444 27804
rect 17948 27748 18004 27758
rect 17948 27654 18004 27692
rect 17612 27188 17668 27198
rect 17164 27074 17220 27086
rect 17164 27022 17166 27074
rect 17218 27022 17220 27074
rect 17164 26908 17220 27022
rect 17612 27076 17668 27132
rect 18060 27076 18116 27114
rect 17612 27074 18004 27076
rect 17612 27022 17614 27074
rect 17666 27022 18004 27074
rect 17612 27020 18004 27022
rect 17612 27010 17668 27020
rect 17164 26852 17444 26908
rect 17388 26292 17444 26852
rect 17388 26226 17444 26236
rect 17836 26852 17892 26862
rect 17836 26178 17892 26796
rect 17836 26126 17838 26178
rect 17890 26126 17892 26178
rect 17388 26068 17444 26078
rect 17388 25618 17444 26012
rect 17388 25566 17390 25618
rect 17442 25566 17444 25618
rect 17388 25554 17444 25566
rect 17500 25956 17556 25966
rect 17052 25454 17054 25506
rect 17106 25454 17108 25506
rect 16380 22878 16382 22930
rect 16434 22878 16436 22930
rect 16380 22866 16436 22878
rect 16492 23156 16548 23166
rect 15708 22652 16100 22708
rect 15820 22484 15876 22494
rect 15820 22370 15876 22428
rect 15820 22318 15822 22370
rect 15874 22318 15876 22370
rect 15708 22148 15764 22158
rect 15708 22054 15764 22092
rect 15148 20132 15204 20972
rect 15148 20038 15204 20076
rect 15260 20972 15540 21028
rect 15596 21474 15652 21486
rect 15596 21422 15598 21474
rect 15650 21422 15652 21474
rect 15036 19348 15092 19386
rect 15036 19282 15092 19292
rect 15260 19236 15316 20972
rect 14868 19180 14980 19236
rect 15148 19234 15316 19236
rect 15148 19182 15262 19234
rect 15314 19182 15316 19234
rect 15148 19180 15316 19182
rect 14812 19170 14868 19180
rect 15036 19124 15092 19134
rect 14700 18284 14980 18340
rect 14364 16882 14420 18284
rect 14588 17668 14644 17678
rect 14588 17666 14868 17668
rect 14588 17614 14590 17666
rect 14642 17614 14868 17666
rect 14588 17612 14868 17614
rect 14588 17602 14644 17612
rect 14476 17444 14532 17454
rect 14476 17350 14532 17388
rect 14364 16830 14366 16882
rect 14418 16830 14420 16882
rect 14364 16818 14420 16830
rect 14476 17220 14532 17230
rect 14476 16098 14532 17164
rect 14812 16658 14868 17612
rect 14924 17444 14980 18284
rect 15036 17666 15092 19068
rect 15036 17614 15038 17666
rect 15090 17614 15092 17666
rect 15036 17602 15092 17614
rect 14924 17388 15092 17444
rect 14812 16606 14814 16658
rect 14866 16606 14868 16658
rect 14476 16046 14478 16098
rect 14530 16046 14532 16098
rect 14476 15988 14532 16046
rect 14476 15922 14532 15932
rect 14588 16436 14644 16446
rect 14588 15986 14644 16380
rect 14588 15934 14590 15986
rect 14642 15934 14644 15986
rect 14252 15474 14308 15484
rect 14140 15262 14142 15314
rect 14194 15262 14196 15314
rect 14140 15250 14196 15262
rect 14252 15316 14308 15326
rect 13916 14366 13918 14418
rect 13970 14366 13972 14418
rect 13916 14354 13972 14366
rect 14028 12964 14084 12974
rect 14028 12870 14084 12908
rect 14028 12290 14084 12302
rect 14028 12238 14030 12290
rect 14082 12238 14084 12290
rect 14028 12068 14084 12238
rect 14028 12002 14084 12012
rect 13804 11340 13972 11396
rect 13804 11172 13860 11182
rect 13692 11170 13860 11172
rect 13692 11118 13806 11170
rect 13858 11118 13860 11170
rect 13692 11116 13860 11118
rect 13468 10610 13524 10622
rect 13468 10558 13470 10610
rect 13522 10558 13524 10610
rect 13468 10500 13524 10558
rect 13468 10434 13524 10444
rect 13580 10612 13636 10622
rect 13580 9938 13636 10556
rect 13580 9886 13582 9938
rect 13634 9886 13636 9938
rect 13580 9874 13636 9886
rect 13692 9826 13748 9838
rect 13692 9774 13694 9826
rect 13746 9774 13748 9826
rect 13692 9716 13748 9774
rect 13804 9828 13860 11116
rect 13804 9762 13860 9772
rect 13692 9650 13748 9660
rect 13916 9492 13972 11340
rect 14028 11060 14084 11070
rect 14028 10722 14084 11004
rect 14252 10834 14308 15260
rect 14588 14644 14644 15934
rect 14476 14196 14532 14206
rect 14476 11788 14532 14140
rect 14588 12852 14644 14588
rect 14812 14196 14868 16606
rect 14924 16996 14980 17006
rect 14924 16770 14980 16940
rect 14924 16718 14926 16770
rect 14978 16718 14980 16770
rect 14924 16548 14980 16718
rect 14924 16482 14980 16492
rect 15036 16436 15092 17388
rect 15148 17108 15204 19180
rect 15260 19170 15316 19180
rect 15372 20804 15428 20814
rect 15260 18338 15316 18350
rect 15260 18286 15262 18338
rect 15314 18286 15316 18338
rect 15260 18228 15316 18286
rect 15260 18162 15316 18172
rect 15372 18004 15428 20748
rect 15596 19908 15652 21422
rect 15820 20802 15876 22318
rect 15820 20750 15822 20802
rect 15874 20750 15876 20802
rect 15820 20132 15876 20750
rect 15820 20066 15876 20076
rect 15596 19842 15652 19852
rect 15932 19234 15988 19246
rect 15932 19182 15934 19234
rect 15986 19182 15988 19234
rect 15708 19124 15764 19134
rect 15708 19030 15764 19068
rect 15820 18562 15876 18574
rect 15820 18510 15822 18562
rect 15874 18510 15876 18562
rect 15148 17042 15204 17052
rect 15260 17948 15428 18004
rect 15484 18450 15540 18462
rect 15484 18398 15486 18450
rect 15538 18398 15540 18450
rect 15260 16882 15316 17948
rect 15484 17556 15540 18398
rect 15820 17780 15876 18510
rect 15820 17686 15876 17724
rect 15932 17892 15988 19182
rect 15540 17500 15652 17556
rect 15484 17490 15540 17500
rect 15372 17108 15428 17118
rect 15428 17052 15540 17108
rect 15372 17042 15428 17052
rect 15260 16830 15262 16882
rect 15314 16830 15316 16882
rect 15260 16818 15316 16830
rect 15372 16884 15428 16894
rect 15036 16370 15092 16380
rect 14700 14140 14868 14196
rect 14924 16324 14980 16334
rect 14924 15428 14980 16268
rect 15260 16212 15316 16222
rect 15260 16118 15316 16156
rect 14924 14196 14980 15372
rect 14700 13860 14756 14140
rect 14924 14130 14980 14140
rect 15148 15986 15204 15998
rect 15148 15934 15150 15986
rect 15202 15934 15204 15986
rect 15148 13972 15204 15934
rect 15260 15092 15316 15102
rect 15260 14998 15316 15036
rect 15260 14532 15316 14542
rect 15372 14532 15428 16828
rect 15484 16882 15540 17052
rect 15484 16830 15486 16882
rect 15538 16830 15540 16882
rect 15484 16818 15540 16830
rect 15484 16212 15540 16222
rect 15484 15652 15540 16156
rect 15596 16100 15652 17500
rect 15932 17220 15988 17836
rect 15932 17154 15988 17164
rect 15932 16884 15988 16894
rect 16044 16884 16100 22652
rect 16268 22372 16324 22382
rect 16492 22372 16548 23100
rect 16268 22370 16548 22372
rect 16268 22318 16270 22370
rect 16322 22318 16548 22370
rect 16268 22316 16548 22318
rect 16604 23042 16660 24332
rect 16940 23938 16996 23950
rect 16940 23886 16942 23938
rect 16994 23886 16996 23938
rect 16828 23828 16884 23838
rect 16828 23734 16884 23772
rect 16940 23716 16996 23886
rect 16940 23650 16996 23660
rect 16940 23492 16996 23502
rect 16604 22990 16606 23042
rect 16658 22990 16660 23042
rect 16268 22306 16324 22316
rect 16604 21924 16660 22990
rect 16716 23156 16772 23166
rect 16716 22484 16772 23100
rect 16940 22708 16996 23436
rect 17052 23044 17108 25454
rect 17500 25508 17556 25900
rect 17836 25620 17892 26126
rect 17836 25554 17892 25564
rect 17500 24946 17556 25452
rect 17948 25506 18004 27020
rect 18060 27010 18116 27020
rect 18396 27074 18452 28700
rect 18620 28690 18676 28700
rect 19292 28690 19348 28702
rect 19740 28644 19796 28654
rect 19740 28550 19796 28588
rect 20524 28644 20580 28654
rect 18956 28532 19012 28542
rect 18956 28082 19012 28476
rect 20524 28530 20580 28588
rect 20524 28478 20526 28530
rect 20578 28478 20580 28530
rect 20300 28420 20356 28430
rect 20300 28326 20356 28364
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 18956 28030 18958 28082
rect 19010 28030 19012 28082
rect 18956 28018 19012 28030
rect 18396 27022 18398 27074
rect 18450 27022 18452 27074
rect 18396 26908 18452 27022
rect 18060 26852 18452 26908
rect 18508 27746 18564 27758
rect 18508 27694 18510 27746
rect 18562 27694 18564 27746
rect 18060 26180 18116 26852
rect 18060 26114 18116 26124
rect 18172 26292 18228 26302
rect 18172 25844 18228 26236
rect 18284 26292 18340 26302
rect 18508 26292 18564 27694
rect 19404 27748 19460 27758
rect 18844 26962 18900 26974
rect 18844 26910 18846 26962
rect 18898 26910 18900 26962
rect 18732 26628 18788 26638
rect 18284 26290 18564 26292
rect 18284 26238 18286 26290
rect 18338 26238 18564 26290
rect 18284 26236 18564 26238
rect 18620 26292 18676 26302
rect 18284 26180 18340 26236
rect 18620 26198 18676 26236
rect 18284 26114 18340 26124
rect 18172 25788 18340 25844
rect 17948 25454 17950 25506
rect 18002 25454 18004 25506
rect 17948 25442 18004 25454
rect 18172 25620 18228 25630
rect 17500 24894 17502 24946
rect 17554 24894 17556 24946
rect 17388 24164 17444 24174
rect 17388 23828 17444 24108
rect 17388 23762 17444 23772
rect 17052 22978 17108 22988
rect 17276 23380 17332 23390
rect 17500 23380 17556 24894
rect 17612 25394 17668 25406
rect 17612 25342 17614 25394
rect 17666 25342 17668 25394
rect 17612 24276 17668 25342
rect 17724 25396 17780 25406
rect 17724 25302 17780 25340
rect 17836 25284 17892 25294
rect 17612 24210 17668 24220
rect 17724 24724 17780 24734
rect 17724 23714 17780 24668
rect 17836 24722 17892 25228
rect 17836 24670 17838 24722
rect 17890 24670 17892 24722
rect 17836 24658 17892 24670
rect 17836 24164 17892 24174
rect 17836 23938 17892 24108
rect 18172 24052 18228 25564
rect 18172 23986 18228 23996
rect 17836 23886 17838 23938
rect 17890 23886 17892 23938
rect 17836 23874 17892 23886
rect 17724 23662 17726 23714
rect 17778 23662 17780 23714
rect 17724 23650 17780 23662
rect 17612 23380 17668 23390
rect 17500 23324 17612 23380
rect 17276 22932 17332 23324
rect 17612 23286 17668 23324
rect 18060 23156 18116 23166
rect 18060 23062 18116 23100
rect 17052 22708 17108 22718
rect 16940 22652 17052 22708
rect 16716 22390 16772 22428
rect 16604 21858 16660 21868
rect 16156 21588 16212 21598
rect 16156 21494 16212 21532
rect 16604 21476 16660 21486
rect 16492 21474 16660 21476
rect 16492 21422 16606 21474
rect 16658 21422 16660 21474
rect 16492 21420 16660 21422
rect 16268 20802 16324 20814
rect 16268 20750 16270 20802
rect 16322 20750 16324 20802
rect 16268 20356 16324 20750
rect 16268 20290 16324 20300
rect 16492 20802 16548 21420
rect 16604 21410 16660 21420
rect 16716 21028 16772 21038
rect 16716 20914 16772 20972
rect 17052 21026 17108 22652
rect 17276 22370 17332 22876
rect 18172 22820 18228 22830
rect 17276 22318 17278 22370
rect 17330 22318 17332 22370
rect 17276 22306 17332 22318
rect 17612 22482 17668 22494
rect 17612 22430 17614 22482
rect 17666 22430 17668 22482
rect 17052 20974 17054 21026
rect 17106 20974 17108 21026
rect 17052 20962 17108 20974
rect 17612 21028 17668 22430
rect 18060 22370 18116 22382
rect 18060 22318 18062 22370
rect 18114 22318 18116 22370
rect 17724 21812 17780 21822
rect 18060 21812 18116 22318
rect 18172 22258 18228 22764
rect 18172 22206 18174 22258
rect 18226 22206 18228 22258
rect 18172 22194 18228 22206
rect 17780 21756 18116 21812
rect 17724 21718 17780 21756
rect 18284 21700 18340 25788
rect 18396 25282 18452 25294
rect 18396 25230 18398 25282
rect 18450 25230 18452 25282
rect 18396 24722 18452 25230
rect 18396 24670 18398 24722
rect 18450 24670 18452 24722
rect 18396 24658 18452 24670
rect 18396 24276 18452 24286
rect 18396 23938 18452 24220
rect 18508 24052 18564 24062
rect 18564 23996 18676 24052
rect 18508 23958 18564 23996
rect 18396 23886 18398 23938
rect 18450 23886 18452 23938
rect 18396 23044 18452 23886
rect 18396 22988 18564 23044
rect 18284 21644 18452 21700
rect 18284 21476 18340 21486
rect 18284 21382 18340 21420
rect 18172 21140 18228 21150
rect 17612 20972 17780 21028
rect 16716 20862 16718 20914
rect 16770 20862 16772 20914
rect 16716 20850 16772 20862
rect 16492 20750 16494 20802
rect 16546 20750 16548 20802
rect 16268 19124 16324 19134
rect 16268 19122 16436 19124
rect 16268 19070 16270 19122
rect 16322 19070 16436 19122
rect 16268 19068 16436 19070
rect 16268 19058 16324 19068
rect 16268 18564 16324 18574
rect 16268 18470 16324 18508
rect 16156 17108 16212 17118
rect 16212 17052 16324 17108
rect 16156 17042 16212 17052
rect 16268 16994 16324 17052
rect 16268 16942 16270 16994
rect 16322 16942 16324 16994
rect 16268 16930 16324 16942
rect 15988 16828 16100 16884
rect 15932 16818 15988 16828
rect 15596 16098 16212 16100
rect 15596 16046 15598 16098
rect 15650 16046 16212 16098
rect 15596 16044 16212 16046
rect 15596 16034 15652 16044
rect 15484 15596 15764 15652
rect 15484 15316 15540 15354
rect 15484 15250 15540 15260
rect 15596 15202 15652 15214
rect 15596 15150 15598 15202
rect 15650 15150 15652 15202
rect 15316 14476 15428 14532
rect 15484 14980 15540 14990
rect 15260 14438 15316 14476
rect 15148 13916 15316 13972
rect 14700 13804 14868 13860
rect 14588 12786 14644 12796
rect 14476 11732 14644 11788
rect 14252 10782 14254 10834
rect 14306 10782 14308 10834
rect 14252 10770 14308 10782
rect 14028 10670 14030 10722
rect 14082 10670 14084 10722
rect 14028 10658 14084 10670
rect 13468 9436 13972 9492
rect 14252 9828 14308 9838
rect 13468 9268 13524 9436
rect 13468 9154 13524 9212
rect 13468 9102 13470 9154
rect 13522 9102 13524 9154
rect 13356 8818 13412 8830
rect 13356 8766 13358 8818
rect 13410 8766 13412 8818
rect 13132 8428 13300 8484
rect 12236 7982 12238 8034
rect 12290 7982 12292 8034
rect 12236 7586 12292 7982
rect 12236 7534 12238 7586
rect 12290 7534 12292 7586
rect 12236 7522 12292 7534
rect 12572 8034 12628 8046
rect 12572 7982 12574 8034
rect 12626 7982 12628 8034
rect 12236 7028 12292 7038
rect 12124 6972 12236 7028
rect 11900 6626 11956 6636
rect 12236 6690 12292 6972
rect 12236 6638 12238 6690
rect 12290 6638 12292 6690
rect 12236 6626 12292 6638
rect 11900 6468 11956 6478
rect 11900 6466 12068 6468
rect 11900 6414 11902 6466
rect 11954 6414 12068 6466
rect 11900 6412 12068 6414
rect 11900 6402 11956 6412
rect 11900 5794 11956 5806
rect 11900 5742 11902 5794
rect 11954 5742 11956 5794
rect 11900 5572 11956 5742
rect 11900 5506 11956 5516
rect 12012 3892 12068 6412
rect 12348 6132 12404 6142
rect 12348 6038 12404 6076
rect 12572 5572 12628 7982
rect 12796 6690 12852 6702
rect 12796 6638 12798 6690
rect 12850 6638 12852 6690
rect 12684 6468 12740 6478
rect 12684 6130 12740 6412
rect 12684 6078 12686 6130
rect 12738 6078 12740 6130
rect 12684 6066 12740 6078
rect 12572 5506 12628 5516
rect 12796 5348 12852 6638
rect 13132 5794 13188 5806
rect 13132 5742 13134 5794
rect 13186 5742 13188 5794
rect 13132 5684 13188 5742
rect 12796 5282 12852 5292
rect 13020 5628 13132 5684
rect 13020 5234 13076 5628
rect 13132 5618 13188 5628
rect 13020 5182 13022 5234
rect 13074 5182 13076 5234
rect 13020 5170 13076 5182
rect 12012 3826 12068 3836
rect 11900 2884 11956 2894
rect 11788 2828 11900 2884
rect 11900 2818 11956 2828
rect 13244 2772 13300 8428
rect 13356 8148 13412 8766
rect 13468 8484 13524 9102
rect 13916 9156 13972 9166
rect 13916 8930 13972 9100
rect 13916 8878 13918 8930
rect 13970 8878 13972 8930
rect 13916 8866 13972 8878
rect 13468 8418 13524 8428
rect 14028 8372 14084 8382
rect 13804 8260 13860 8270
rect 13804 8166 13860 8204
rect 13356 8082 13412 8092
rect 13468 7476 13524 7486
rect 13468 7382 13524 7420
rect 13580 7364 13636 7374
rect 13468 6804 13524 6814
rect 13580 6804 13636 7308
rect 14028 6916 14084 8316
rect 14252 6916 14308 9772
rect 14476 9714 14532 9726
rect 14476 9662 14478 9714
rect 14530 9662 14532 9714
rect 14476 9380 14532 9662
rect 14476 9314 14532 9324
rect 14364 9268 14420 9278
rect 14364 9174 14420 9212
rect 14364 8260 14420 8270
rect 14364 8166 14420 8204
rect 14588 7588 14644 11732
rect 14700 9940 14756 9950
rect 14700 9846 14756 9884
rect 14812 9716 14868 13804
rect 14924 13748 14980 13786
rect 14924 13682 14980 13692
rect 15036 13188 15092 13198
rect 15036 11506 15092 13132
rect 15148 13188 15204 13226
rect 15148 13122 15204 13132
rect 15260 12740 15316 13916
rect 15036 11454 15038 11506
rect 15090 11454 15092 11506
rect 15036 11442 15092 11454
rect 15148 12684 15316 12740
rect 15484 13746 15540 14924
rect 15484 13694 15486 13746
rect 15538 13694 15540 13746
rect 15148 10610 15204 12684
rect 15372 12516 15428 12526
rect 15260 12404 15316 12414
rect 15260 12178 15316 12348
rect 15260 12126 15262 12178
rect 15314 12126 15316 12178
rect 15260 12114 15316 12126
rect 15148 10558 15150 10610
rect 15202 10558 15204 10610
rect 15148 10546 15204 10558
rect 15260 11394 15316 11406
rect 15260 11342 15262 11394
rect 15314 11342 15316 11394
rect 15260 10164 15316 11342
rect 15372 10610 15428 12460
rect 15484 12402 15540 13694
rect 15596 13188 15652 15150
rect 15596 13122 15652 13132
rect 15484 12350 15486 12402
rect 15538 12350 15540 12402
rect 15484 12338 15540 12350
rect 15372 10558 15374 10610
rect 15426 10558 15428 10610
rect 15372 10546 15428 10558
rect 15484 11844 15540 11854
rect 15036 10108 15316 10164
rect 15372 10388 15428 10398
rect 14588 7494 14644 7532
rect 14700 9660 14868 9716
rect 14924 10052 14980 10062
rect 14924 9826 14980 9996
rect 14924 9774 14926 9826
rect 14978 9774 14980 9826
rect 14252 6860 14420 6916
rect 14028 6822 14084 6860
rect 13524 6748 13636 6804
rect 13468 6738 13524 6748
rect 13468 5682 13524 5694
rect 13468 5630 13470 5682
rect 13522 5630 13524 5682
rect 13468 5572 13524 5630
rect 13468 5506 13524 5516
rect 13580 5236 13636 6748
rect 13692 6692 13748 6702
rect 13692 6130 13748 6636
rect 13692 6078 13694 6130
rect 13746 6078 13748 6130
rect 13692 6066 13748 6078
rect 13804 6690 13860 6702
rect 13804 6638 13806 6690
rect 13858 6638 13860 6690
rect 13804 5794 13860 6638
rect 14252 6690 14308 6702
rect 14252 6638 14254 6690
rect 14306 6638 14308 6690
rect 14252 6130 14308 6638
rect 14252 6078 14254 6130
rect 14306 6078 14308 6130
rect 14252 6066 14308 6078
rect 13804 5742 13806 5794
rect 13858 5742 13860 5794
rect 13804 5730 13860 5742
rect 14364 5460 14420 6860
rect 14700 6914 14756 9660
rect 14812 9380 14868 9390
rect 14812 9042 14868 9324
rect 14924 9156 14980 9774
rect 14924 9062 14980 9100
rect 14812 8990 14814 9042
rect 14866 8990 14868 9042
rect 14812 8978 14868 8990
rect 14812 8484 14868 8494
rect 15036 8484 15092 10108
rect 15372 10052 15428 10332
rect 14812 8482 15092 8484
rect 14812 8430 14814 8482
rect 14866 8430 15092 8482
rect 14812 8428 15092 8430
rect 15260 9996 15428 10052
rect 14812 8418 14868 8428
rect 14924 8258 14980 8270
rect 14924 8206 14926 8258
rect 14978 8206 14980 8258
rect 14924 8036 14980 8206
rect 15260 8258 15316 9996
rect 15484 9828 15540 11788
rect 15708 11620 15764 15596
rect 15260 8206 15262 8258
rect 15314 8206 15316 8258
rect 15260 8194 15316 8206
rect 15372 9772 15540 9828
rect 15596 10724 15652 10734
rect 15596 10610 15652 10668
rect 15596 10558 15598 10610
rect 15650 10558 15652 10610
rect 15372 8260 15428 9772
rect 15372 8194 15428 8204
rect 15484 9602 15540 9614
rect 15484 9550 15486 9602
rect 15538 9550 15540 9602
rect 15484 9268 15540 9550
rect 15372 8036 15428 8046
rect 14924 7980 15316 8036
rect 15260 7924 15316 7980
rect 15260 7252 15316 7868
rect 15372 7698 15428 7980
rect 15372 7646 15374 7698
rect 15426 7646 15428 7698
rect 15372 7634 15428 7646
rect 15484 7700 15540 9212
rect 15596 8708 15652 10558
rect 15708 10388 15764 11564
rect 15932 14420 15988 14430
rect 15932 12628 15988 14364
rect 15708 10322 15764 10332
rect 15820 11284 15876 11294
rect 15820 9826 15876 11228
rect 15820 9774 15822 9826
rect 15874 9774 15876 9826
rect 15820 9762 15876 9774
rect 15932 9604 15988 12572
rect 16044 13522 16100 13534
rect 16044 13470 16046 13522
rect 16098 13470 16100 13522
rect 16044 11394 16100 13470
rect 16156 12964 16212 16044
rect 16380 14084 16436 19068
rect 16492 17332 16548 20750
rect 17388 20802 17444 20814
rect 17388 20750 17390 20802
rect 17442 20750 17444 20802
rect 16604 20692 16660 20702
rect 16604 20242 16660 20636
rect 16828 20690 16884 20702
rect 16828 20638 16830 20690
rect 16882 20638 16884 20690
rect 16604 20190 16606 20242
rect 16658 20190 16660 20242
rect 16604 20178 16660 20190
rect 16716 20580 16772 20590
rect 16604 20018 16660 20030
rect 16604 19966 16606 20018
rect 16658 19966 16660 20018
rect 16604 19684 16660 19966
rect 16716 20020 16772 20524
rect 16716 19954 16772 19964
rect 16604 19460 16660 19628
rect 16604 19394 16660 19404
rect 16604 19012 16660 19022
rect 16604 18116 16660 18956
rect 16828 18676 16884 20638
rect 17388 20356 17444 20750
rect 17612 20804 17668 20814
rect 17612 20710 17668 20748
rect 17724 20468 17780 20972
rect 18172 20914 18228 21084
rect 18172 20862 18174 20914
rect 18226 20862 18228 20914
rect 18172 20850 18228 20862
rect 17724 20402 17780 20412
rect 17948 20804 18004 20814
rect 17388 20290 17444 20300
rect 17836 20356 17892 20366
rect 16940 20020 16996 20030
rect 16940 19122 16996 19964
rect 17612 20020 17668 20030
rect 17612 19908 17668 19964
rect 17612 19906 17780 19908
rect 17612 19854 17614 19906
rect 17666 19854 17780 19906
rect 17612 19852 17780 19854
rect 17612 19842 17668 19852
rect 17500 19796 17556 19806
rect 16940 19070 16942 19122
rect 16994 19070 16996 19122
rect 16940 19058 16996 19070
rect 17164 19460 17220 19470
rect 17164 19124 17220 19404
rect 17500 19458 17556 19740
rect 17500 19406 17502 19458
rect 17554 19406 17556 19458
rect 17164 19058 17220 19068
rect 17276 19122 17332 19134
rect 17276 19070 17278 19122
rect 17330 19070 17332 19122
rect 16716 18564 16772 18574
rect 16716 18470 16772 18508
rect 16604 18050 16660 18060
rect 16828 17554 16884 18620
rect 17276 18340 17332 19070
rect 17500 19124 17556 19406
rect 17500 19058 17556 19068
rect 16940 18116 16996 18126
rect 16940 17668 16996 18060
rect 16940 17602 16996 17612
rect 16828 17502 16830 17554
rect 16882 17502 16884 17554
rect 16828 17490 16884 17502
rect 17052 17554 17108 17566
rect 17052 17502 17054 17554
rect 17106 17502 17108 17554
rect 17052 17444 17108 17502
rect 17276 17556 17332 18284
rect 17612 18562 17668 18574
rect 17612 18510 17614 18562
rect 17666 18510 17668 18562
rect 17612 18452 17668 18510
rect 17724 18564 17780 19852
rect 17836 19458 17892 20300
rect 17948 19908 18004 20748
rect 18060 20132 18116 20142
rect 18060 20038 18116 20076
rect 17948 19852 18116 19908
rect 17836 19406 17838 19458
rect 17890 19406 17892 19458
rect 17836 19394 17892 19406
rect 17724 18508 17892 18564
rect 17276 17490 17332 17500
rect 17388 18226 17444 18238
rect 17388 18174 17390 18226
rect 17442 18174 17444 18226
rect 16940 17388 17108 17444
rect 16604 17332 16660 17342
rect 16492 17276 16604 17332
rect 16492 16212 16548 16222
rect 16492 16118 16548 16156
rect 16604 14530 16660 17276
rect 16828 16884 16884 16894
rect 16828 16790 16884 16828
rect 16828 16548 16884 16558
rect 16828 16098 16884 16492
rect 16940 16324 16996 17388
rect 17388 17332 17444 18174
rect 17612 18004 17668 18396
rect 17724 18340 17780 18350
rect 17724 18246 17780 18284
rect 17612 17938 17668 17948
rect 17388 17266 17444 17276
rect 17612 17666 17668 17678
rect 17612 17614 17614 17666
rect 17666 17614 17668 17666
rect 17612 17220 17668 17614
rect 17724 17668 17780 17678
rect 17724 17574 17780 17612
rect 17612 17154 17668 17164
rect 17724 17444 17780 17454
rect 17724 16994 17780 17388
rect 17724 16942 17726 16994
rect 17778 16942 17780 16994
rect 17724 16930 17780 16942
rect 17500 16436 17556 16446
rect 16940 16268 17108 16324
rect 16828 16046 16830 16098
rect 16882 16046 16884 16098
rect 16828 16034 16884 16046
rect 16940 16100 16996 16110
rect 16940 15876 16996 16044
rect 16940 15652 16996 15820
rect 16604 14478 16606 14530
rect 16658 14478 16660 14530
rect 16604 14466 16660 14478
rect 16828 15596 16996 15652
rect 16380 14028 16660 14084
rect 16268 13748 16324 13758
rect 16268 13654 16324 13692
rect 16604 13076 16660 14028
rect 16604 13074 16772 13076
rect 16604 13022 16606 13074
rect 16658 13022 16772 13074
rect 16604 13020 16772 13022
rect 16604 13010 16660 13020
rect 16268 12964 16324 12974
rect 16156 12962 16324 12964
rect 16156 12910 16270 12962
rect 16322 12910 16324 12962
rect 16156 12908 16324 12910
rect 16268 12898 16324 12908
rect 16604 12740 16660 12750
rect 16492 12684 16604 12740
rect 16380 12516 16436 12526
rect 16044 11342 16046 11394
rect 16098 11342 16100 11394
rect 16044 11330 16100 11342
rect 16156 11732 16212 11742
rect 16156 10612 16212 11676
rect 16380 10834 16436 12460
rect 16380 10782 16382 10834
rect 16434 10782 16436 10834
rect 16380 10770 16436 10782
rect 15988 9548 16100 9604
rect 15932 9538 15988 9548
rect 15596 8642 15652 8652
rect 15708 9380 15764 9390
rect 15708 8596 15764 9324
rect 15820 9268 15876 9278
rect 15820 9174 15876 9212
rect 15932 9156 15988 9166
rect 16044 9156 16100 9548
rect 16156 9268 16212 10556
rect 16268 9268 16324 9278
rect 16156 9266 16324 9268
rect 16156 9214 16270 9266
rect 16322 9214 16324 9266
rect 16156 9212 16324 9214
rect 16268 9202 16324 9212
rect 16380 9268 16436 9278
rect 16492 9268 16548 12684
rect 16604 12674 16660 12684
rect 16716 11956 16772 13020
rect 16716 11890 16772 11900
rect 16828 12402 16884 15596
rect 16940 15428 16996 15438
rect 16940 13970 16996 15372
rect 16940 13918 16942 13970
rect 16994 13918 16996 13970
rect 16940 13906 16996 13918
rect 16828 12350 16830 12402
rect 16882 12350 16884 12402
rect 16716 11732 16772 11742
rect 16716 11284 16772 11676
rect 16380 9266 16548 9268
rect 16380 9214 16382 9266
rect 16434 9214 16548 9266
rect 16380 9212 16548 9214
rect 16604 11228 16716 11284
rect 16380 9202 16436 9212
rect 16044 9100 16212 9156
rect 15932 9042 15988 9100
rect 15932 8990 15934 9042
rect 15986 8990 15988 9042
rect 15932 8978 15988 8990
rect 16156 9044 16212 9100
rect 16492 9044 16548 9054
rect 16212 9042 16548 9044
rect 16212 8990 16494 9042
rect 16546 8990 16548 9042
rect 16212 8988 16548 8990
rect 16156 8950 16212 8988
rect 16492 8978 16548 8988
rect 15708 8530 15764 8540
rect 15820 8820 15876 8830
rect 15484 7634 15540 7644
rect 15484 7476 15540 7486
rect 15484 7382 15540 7420
rect 15260 7196 15652 7252
rect 14700 6862 14702 6914
rect 14754 6862 14756 6914
rect 14700 6850 14756 6862
rect 14476 6804 14532 6814
rect 14476 6132 14532 6748
rect 15036 6690 15092 6702
rect 15036 6638 15038 6690
rect 15090 6638 15092 6690
rect 14476 6066 14532 6076
rect 14700 6580 14756 6590
rect 14588 5684 14644 5694
rect 14588 5590 14644 5628
rect 14364 5404 14644 5460
rect 13692 5236 13748 5246
rect 13580 5234 13748 5236
rect 13580 5182 13694 5234
rect 13746 5182 13748 5234
rect 13580 5180 13748 5182
rect 13692 5170 13748 5180
rect 14028 5236 14084 5246
rect 14028 5142 14084 5180
rect 14588 5234 14644 5404
rect 14588 5182 14590 5234
rect 14642 5182 14644 5234
rect 14588 5170 14644 5182
rect 14700 5124 14756 6524
rect 14812 5796 14868 5806
rect 14812 5794 14980 5796
rect 14812 5742 14814 5794
rect 14866 5742 14980 5794
rect 14812 5740 14980 5742
rect 14812 5730 14868 5740
rect 14812 5348 14868 5358
rect 14812 5254 14868 5292
rect 14924 5124 14980 5740
rect 15036 5348 15092 6638
rect 15148 6466 15204 6478
rect 15484 6468 15540 6478
rect 15148 6414 15150 6466
rect 15202 6414 15204 6466
rect 15148 6020 15204 6414
rect 15148 5954 15204 5964
rect 15260 6466 15540 6468
rect 15260 6414 15486 6466
rect 15538 6414 15540 6466
rect 15260 6412 15540 6414
rect 15260 6018 15316 6412
rect 15484 6402 15540 6412
rect 15596 6244 15652 7196
rect 15820 6690 15876 8764
rect 16492 8596 16548 8606
rect 15932 8372 15988 8382
rect 15932 8258 15988 8316
rect 16380 8372 16436 8382
rect 15932 8206 15934 8258
rect 15986 8206 15988 8258
rect 15932 8194 15988 8206
rect 16268 8260 16324 8270
rect 16268 8166 16324 8204
rect 16156 8148 16212 8158
rect 16044 8092 16156 8148
rect 16044 8034 16100 8092
rect 16156 8082 16212 8092
rect 16044 7982 16046 8034
rect 16098 7982 16100 8034
rect 16044 7970 16100 7982
rect 15932 7700 15988 7710
rect 15932 7474 15988 7644
rect 16380 7586 16436 8316
rect 16380 7534 16382 7586
rect 16434 7534 16436 7586
rect 16380 7522 16436 7534
rect 15932 7422 15934 7474
rect 15986 7422 15988 7474
rect 15932 7410 15988 7422
rect 16044 7474 16100 7486
rect 16044 7422 16046 7474
rect 16098 7422 16100 7474
rect 15820 6638 15822 6690
rect 15874 6638 15876 6690
rect 15260 5966 15262 6018
rect 15314 5966 15316 6018
rect 15260 5954 15316 5966
rect 15484 6188 15652 6244
rect 15708 6580 15764 6590
rect 15708 6466 15764 6524
rect 15708 6414 15710 6466
rect 15762 6414 15764 6466
rect 15484 5906 15540 6188
rect 15484 5854 15486 5906
rect 15538 5854 15540 5906
rect 15484 5842 15540 5854
rect 15596 5908 15652 5918
rect 15484 5348 15540 5358
rect 15036 5346 15540 5348
rect 15036 5294 15486 5346
rect 15538 5294 15540 5346
rect 15036 5292 15540 5294
rect 15484 5282 15540 5292
rect 14700 5068 14868 5124
rect 14924 5068 15092 5124
rect 14364 5012 14420 5022
rect 14364 4562 14420 4956
rect 14364 4510 14366 4562
rect 14418 4510 14420 4562
rect 14364 4498 14420 4510
rect 14700 4226 14756 4238
rect 14700 4174 14702 4226
rect 14754 4174 14756 4226
rect 14700 3892 14756 4174
rect 14700 3826 14756 3836
rect 14812 3668 14868 5068
rect 15036 5012 15092 5068
rect 15148 5122 15204 5134
rect 15148 5070 15150 5122
rect 15202 5070 15204 5122
rect 15148 5012 15204 5070
rect 15260 5124 15316 5134
rect 15260 5012 15316 5068
rect 15484 5124 15540 5134
rect 15596 5124 15652 5852
rect 15708 5796 15764 6414
rect 15820 6468 15876 6638
rect 15820 6402 15876 6412
rect 16044 6692 16100 7422
rect 16156 7476 16212 7486
rect 16156 6802 16212 7420
rect 16268 7364 16324 7374
rect 16268 7270 16324 7308
rect 16492 6916 16548 8540
rect 16604 8036 16660 11228
rect 16716 11218 16772 11228
rect 16828 10836 16884 12350
rect 16940 13636 16996 13646
rect 16940 11844 16996 13580
rect 17052 12404 17108 16268
rect 17164 16212 17220 16222
rect 17164 16118 17220 16156
rect 17500 15540 17556 16380
rect 17836 16100 17892 18508
rect 17948 17666 18004 17678
rect 17948 17614 17950 17666
rect 18002 17614 18004 17666
rect 17948 17332 18004 17614
rect 17948 17266 18004 17276
rect 17948 17108 18004 17118
rect 17948 16994 18004 17052
rect 17948 16942 17950 16994
rect 18002 16942 18004 16994
rect 17948 16884 18004 16942
rect 17948 16818 18004 16828
rect 17948 16548 18004 16558
rect 18060 16548 18116 19852
rect 18396 19460 18452 21644
rect 18508 21252 18564 22988
rect 18620 22036 18676 23996
rect 18620 21970 18676 21980
rect 18620 21588 18676 21598
rect 18620 21494 18676 21532
rect 18508 21196 18676 21252
rect 18620 20580 18676 21196
rect 18732 20804 18788 26572
rect 18844 26292 18900 26910
rect 19404 26850 19460 27692
rect 19404 26798 19406 26850
rect 19458 26798 19460 26850
rect 19404 26740 19460 26798
rect 19404 26674 19460 26684
rect 19516 27746 19572 27758
rect 19852 27748 19908 27758
rect 19516 27694 19518 27746
rect 19570 27694 19572 27746
rect 19516 26516 19572 27694
rect 19628 27746 19908 27748
rect 19628 27694 19854 27746
rect 19906 27694 19908 27746
rect 19628 27692 19908 27694
rect 19628 26740 19684 27692
rect 19852 27682 19908 27692
rect 19852 27412 19908 27422
rect 19852 27186 19908 27356
rect 19852 27134 19854 27186
rect 19906 27134 19908 27186
rect 19852 27122 19908 27134
rect 20412 26962 20468 26974
rect 20412 26910 20414 26962
rect 20466 26910 20468 26962
rect 19628 26674 19684 26684
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19516 26460 19908 26516
rect 19852 26404 19908 26460
rect 18844 26226 18900 26236
rect 19068 26290 19124 26302
rect 19068 26238 19070 26290
rect 19122 26238 19124 26290
rect 19068 26180 19124 26238
rect 19740 26292 19796 26302
rect 18956 25282 19012 25294
rect 18956 25230 18958 25282
rect 19010 25230 19012 25282
rect 18956 24500 19012 25230
rect 18956 24434 19012 24444
rect 18844 23266 18900 23278
rect 18844 23214 18846 23266
rect 18898 23214 18900 23266
rect 18844 21812 18900 23214
rect 19068 22372 19124 26124
rect 19404 26180 19460 26190
rect 19404 26178 19572 26180
rect 19404 26126 19406 26178
rect 19458 26126 19572 26178
rect 19404 26124 19572 26126
rect 19404 26114 19460 26124
rect 19516 25620 19572 26124
rect 19516 25554 19572 25564
rect 19740 26178 19796 26236
rect 19740 26126 19742 26178
rect 19794 26126 19796 26178
rect 19292 25396 19348 25406
rect 19740 25396 19796 26126
rect 19852 25732 19908 26348
rect 20188 26292 20244 26302
rect 20188 26198 20244 26236
rect 20412 26180 20468 26910
rect 20524 26908 20580 28478
rect 20636 28530 20692 29596
rect 21196 29652 21252 29662
rect 21196 29426 21252 29596
rect 21196 29374 21198 29426
rect 21250 29374 21252 29426
rect 21196 29362 21252 29374
rect 20748 29316 20804 29326
rect 20748 29222 20804 29260
rect 21308 29316 21364 29326
rect 21308 28642 21364 29260
rect 21420 28754 21476 29932
rect 21532 29922 21588 29932
rect 21756 29988 21812 29998
rect 21756 29894 21812 29932
rect 21980 29652 22036 29662
rect 21980 29558 22036 29596
rect 21644 29426 21700 29438
rect 21644 29374 21646 29426
rect 21698 29374 21700 29426
rect 21644 29316 21700 29374
rect 21644 29250 21700 29260
rect 22092 29204 22148 30156
rect 22204 29540 22260 29550
rect 22204 29446 22260 29484
rect 22316 29540 22372 30156
rect 23772 30212 23828 30222
rect 23772 30118 23828 30156
rect 22540 29988 22596 29998
rect 22316 29538 22484 29540
rect 22316 29486 22318 29538
rect 22370 29486 22484 29538
rect 22316 29484 22484 29486
rect 22316 29474 22372 29484
rect 22316 29204 22372 29214
rect 22092 29202 22372 29204
rect 22092 29150 22318 29202
rect 22370 29150 22372 29202
rect 22092 29148 22372 29150
rect 22316 29138 22372 29148
rect 21420 28702 21422 28754
rect 21474 28702 21476 28754
rect 21420 28690 21476 28702
rect 21980 28756 22036 28766
rect 21308 28590 21310 28642
rect 21362 28590 21364 28642
rect 21308 28578 21364 28590
rect 21644 28644 21700 28654
rect 20636 28478 20638 28530
rect 20690 28478 20692 28530
rect 20636 28466 20692 28478
rect 20860 28418 20916 28430
rect 20860 28366 20862 28418
rect 20914 28366 20916 28418
rect 20524 26852 20692 26908
rect 20524 26404 20580 26414
rect 20524 26310 20580 26348
rect 20412 26114 20468 26124
rect 19852 25666 19908 25676
rect 20188 25508 20244 25518
rect 20188 25414 20244 25452
rect 19180 25394 19348 25396
rect 19180 25342 19294 25394
rect 19346 25342 19348 25394
rect 19180 25340 19348 25342
rect 19180 22596 19236 25340
rect 19292 25330 19348 25340
rect 19516 25340 19796 25396
rect 19404 24836 19460 24846
rect 19404 24162 19460 24780
rect 19404 24110 19406 24162
rect 19458 24110 19460 24162
rect 19404 24098 19460 24110
rect 19292 24050 19348 24062
rect 19292 23998 19294 24050
rect 19346 23998 19348 24050
rect 19292 22820 19348 23998
rect 19404 23938 19460 23950
rect 19404 23886 19406 23938
rect 19458 23886 19460 23938
rect 19404 23828 19460 23886
rect 19404 23762 19460 23772
rect 19516 23380 19572 25340
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20188 24724 20244 24734
rect 20188 24630 20244 24668
rect 19292 22754 19348 22764
rect 19404 23324 19572 23380
rect 19628 24164 19684 24174
rect 19180 22540 19348 22596
rect 19180 22372 19236 22410
rect 19068 22316 19180 22372
rect 19180 22306 19236 22316
rect 18956 22260 19012 22270
rect 18956 22146 19012 22204
rect 18956 22094 18958 22146
rect 19010 22094 19012 22146
rect 18956 22082 19012 22094
rect 18844 21756 19236 21812
rect 18844 21588 18900 21598
rect 18844 21364 18900 21532
rect 18844 21298 18900 21308
rect 19068 21586 19124 21598
rect 19068 21534 19070 21586
rect 19122 21534 19124 21586
rect 19068 21476 19124 21534
rect 18732 20738 18788 20748
rect 18956 21252 19012 21262
rect 18620 20578 18788 20580
rect 18620 20526 18622 20578
rect 18674 20526 18788 20578
rect 18620 20524 18788 20526
rect 18620 20514 18676 20524
rect 18620 20020 18676 20030
rect 18620 19926 18676 19964
rect 18732 19796 18788 20524
rect 18396 19346 18452 19404
rect 18396 19294 18398 19346
rect 18450 19294 18452 19346
rect 18172 17666 18228 17678
rect 18172 17614 18174 17666
rect 18226 17614 18228 17666
rect 18172 16996 18228 17614
rect 18172 16930 18228 16940
rect 18004 16492 18116 16548
rect 17948 16482 18004 16492
rect 17052 12338 17108 12348
rect 17276 15538 17556 15540
rect 17276 15486 17502 15538
rect 17554 15486 17556 15538
rect 17276 15484 17556 15486
rect 17164 11844 17220 11854
rect 16940 11788 17164 11844
rect 16940 11508 16996 11788
rect 17164 11778 17220 11788
rect 16940 11060 16996 11452
rect 16940 10994 16996 11004
rect 17052 11394 17108 11406
rect 17052 11342 17054 11394
rect 17106 11342 17108 11394
rect 16828 10770 16884 10780
rect 16940 10724 16996 10734
rect 16828 10612 16884 10622
rect 16940 10612 16996 10668
rect 16828 10610 16996 10612
rect 16828 10558 16830 10610
rect 16882 10558 16996 10610
rect 16828 10556 16996 10558
rect 16828 10546 16884 10556
rect 17052 10164 17108 11342
rect 16940 10108 17108 10164
rect 17164 11284 17220 11294
rect 16828 9826 16884 9838
rect 16828 9774 16830 9826
rect 16882 9774 16884 9826
rect 16716 9714 16772 9726
rect 16716 9662 16718 9714
rect 16770 9662 16772 9714
rect 16716 9492 16772 9662
rect 16716 9426 16772 9436
rect 16828 9268 16884 9774
rect 16716 9212 16884 9268
rect 16940 9268 16996 10108
rect 17052 9938 17108 9950
rect 17052 9886 17054 9938
rect 17106 9886 17108 9938
rect 17052 9828 17108 9886
rect 17052 9762 17108 9772
rect 16716 8372 16772 9212
rect 16940 9202 16996 9212
rect 17164 9156 17220 11228
rect 17276 10052 17332 15484
rect 17500 15474 17556 15484
rect 17612 16098 17892 16100
rect 17612 16046 17838 16098
rect 17890 16046 17892 16098
rect 17612 16044 17892 16046
rect 17500 14644 17556 14654
rect 17500 14530 17556 14588
rect 17500 14478 17502 14530
rect 17554 14478 17556 14530
rect 17500 14466 17556 14478
rect 17612 13746 17668 16044
rect 17836 16034 17892 16044
rect 18060 16212 18116 16222
rect 17948 15316 18004 15326
rect 17836 14308 17892 14318
rect 17612 13694 17614 13746
rect 17666 13694 17668 13746
rect 17612 13682 17668 13694
rect 17724 14306 17892 14308
rect 17724 14254 17838 14306
rect 17890 14254 17892 14306
rect 17724 14252 17892 14254
rect 17724 13300 17780 14252
rect 17836 14242 17892 14252
rect 17388 13244 17780 13300
rect 17388 12850 17444 13244
rect 17836 13188 17892 13198
rect 17948 13188 18004 15260
rect 18060 14532 18116 16156
rect 18172 15540 18228 15550
rect 18172 15314 18228 15484
rect 18172 15262 18174 15314
rect 18226 15262 18228 15314
rect 18172 15250 18228 15262
rect 18172 14532 18228 14542
rect 18060 14530 18228 14532
rect 18060 14478 18174 14530
rect 18226 14478 18228 14530
rect 18060 14476 18228 14478
rect 18172 14466 18228 14476
rect 18396 14196 18452 19294
rect 18620 19740 18788 19796
rect 18844 20468 18900 20478
rect 18844 19796 18900 20412
rect 18956 20242 19012 21196
rect 18956 20190 18958 20242
rect 19010 20190 19012 20242
rect 18956 20178 19012 20190
rect 18956 19796 19012 19806
rect 18844 19794 19012 19796
rect 18844 19742 18958 19794
rect 19010 19742 19012 19794
rect 18844 19740 19012 19742
rect 18620 19012 18676 19740
rect 18620 18946 18676 18956
rect 18732 19236 18788 19246
rect 18620 18562 18676 18574
rect 18620 18510 18622 18562
rect 18674 18510 18676 18562
rect 18620 18452 18676 18510
rect 18620 17892 18676 18396
rect 18732 18450 18788 19180
rect 18844 19010 18900 19022
rect 18844 18958 18846 19010
rect 18898 18958 18900 19010
rect 18844 18564 18900 18958
rect 18844 18498 18900 18508
rect 18732 18398 18734 18450
rect 18786 18398 18788 18450
rect 18732 18386 18788 18398
rect 18732 17892 18788 17902
rect 18620 17836 18732 17892
rect 18732 17826 18788 17836
rect 18732 17554 18788 17566
rect 18732 17502 18734 17554
rect 18786 17502 18788 17554
rect 18620 17444 18676 17454
rect 18508 17220 18564 17230
rect 18508 16882 18564 17164
rect 18620 16994 18676 17388
rect 18620 16942 18622 16994
rect 18674 16942 18676 16994
rect 18620 16930 18676 16942
rect 18508 16830 18510 16882
rect 18562 16830 18564 16882
rect 18508 14420 18564 16830
rect 18732 15316 18788 17502
rect 18956 17332 19012 19740
rect 19068 19236 19124 21420
rect 19180 20468 19236 21756
rect 19292 21476 19348 22540
rect 19404 22148 19460 23324
rect 19628 23154 19684 24108
rect 20636 24052 20692 26852
rect 20748 26852 20804 26862
rect 20748 26758 20804 26796
rect 20860 26404 20916 28366
rect 21532 28420 21588 28430
rect 21532 28326 21588 28364
rect 21532 27412 21588 27422
rect 21308 26964 21364 27002
rect 21308 26898 21364 26908
rect 20860 26338 20916 26348
rect 21532 26292 21588 27356
rect 21196 26290 21588 26292
rect 21196 26238 21534 26290
rect 21586 26238 21588 26290
rect 21196 26236 21588 26238
rect 20860 26178 20916 26190
rect 20860 26126 20862 26178
rect 20914 26126 20916 26178
rect 20860 25732 20916 26126
rect 20860 25666 20916 25676
rect 21196 25396 21252 26236
rect 21532 26226 21588 26236
rect 20860 25340 21252 25396
rect 21532 25396 21588 25406
rect 21644 25396 21700 28588
rect 21980 28642 22036 28700
rect 21980 28590 21982 28642
rect 22034 28590 22036 28642
rect 21980 28578 22036 28590
rect 22316 28644 22372 28654
rect 22428 28644 22484 29484
rect 22316 28642 22484 28644
rect 22316 28590 22318 28642
rect 22370 28590 22484 28642
rect 22316 28588 22484 28590
rect 22316 28420 22372 28588
rect 22316 28354 22372 28364
rect 22316 27972 22372 27982
rect 21756 27186 21812 27198
rect 21756 27134 21758 27186
rect 21810 27134 21812 27186
rect 21756 26908 21812 27134
rect 22316 27188 22372 27916
rect 22540 27860 22596 29932
rect 23996 29652 24052 30270
rect 23996 29586 24052 29596
rect 22876 29316 22932 29326
rect 22764 28644 22820 28654
rect 22876 28644 22932 29260
rect 24108 28756 24164 30716
rect 24220 30210 24276 32284
rect 24444 31778 24500 31790
rect 24444 31726 24446 31778
rect 24498 31726 24500 31778
rect 24444 30884 24500 31726
rect 24444 30818 24500 30828
rect 25004 31780 25060 31790
rect 25228 31780 25284 31790
rect 25004 31778 25228 31780
rect 25004 31726 25006 31778
rect 25058 31726 25228 31778
rect 25004 31724 25228 31726
rect 24220 30158 24222 30210
rect 24274 30158 24276 30210
rect 24220 30146 24276 30158
rect 24668 30212 24724 30222
rect 24332 29988 24388 29998
rect 24332 29894 24388 29932
rect 24444 29986 24500 29998
rect 24444 29934 24446 29986
rect 24498 29934 24500 29986
rect 24220 29314 24276 29326
rect 24220 29262 24222 29314
rect 24274 29262 24276 29314
rect 24220 29202 24276 29262
rect 24220 29150 24222 29202
rect 24274 29150 24276 29202
rect 24220 29138 24276 29150
rect 24444 29202 24500 29934
rect 24668 29650 24724 30156
rect 25004 30210 25060 31724
rect 25228 31714 25284 31724
rect 25788 31556 25844 31566
rect 25788 31220 25844 31500
rect 25788 31126 25844 31164
rect 25900 31554 25956 32508
rect 26124 32562 26180 32574
rect 26124 32510 26126 32562
rect 26178 32510 26180 32562
rect 26124 31780 26180 32510
rect 26348 32564 26404 33518
rect 26460 33570 26516 33740
rect 26460 33518 26462 33570
rect 26514 33518 26516 33570
rect 26460 33506 26516 33518
rect 26572 33348 26628 33852
rect 27580 33458 27636 34748
rect 28028 33572 28084 36876
rect 28364 36820 28420 38612
rect 28476 38612 28756 38668
rect 28476 37492 28532 38612
rect 29036 38500 29092 40908
rect 29148 40292 29204 42030
rect 29260 42642 29428 42644
rect 29260 42590 29374 42642
rect 29426 42590 29428 42642
rect 29260 42588 29428 42590
rect 29260 41858 29316 42588
rect 29372 42578 29428 42588
rect 29372 41972 29428 41982
rect 29372 41878 29428 41916
rect 29260 41806 29262 41858
rect 29314 41806 29316 41858
rect 29260 41794 29316 41806
rect 29148 40226 29204 40236
rect 29372 39844 29428 39854
rect 29484 39844 29540 44268
rect 29708 44324 29764 44334
rect 29708 44230 29764 44268
rect 29820 44212 29876 44222
rect 29820 44118 29876 44156
rect 29932 43988 29988 45388
rect 29820 43932 29988 43988
rect 30044 44546 30100 45612
rect 30044 44494 30046 44546
rect 30098 44494 30100 44546
rect 29596 43540 29652 43550
rect 29820 43540 29876 43932
rect 29932 43764 29988 43774
rect 29932 43670 29988 43708
rect 30044 43652 30100 44494
rect 30156 45220 30212 45838
rect 30156 43764 30212 45164
rect 30156 43698 30212 43708
rect 30044 43586 30100 43596
rect 29820 43484 29988 43540
rect 29596 43446 29652 43484
rect 29708 43092 29764 43102
rect 29764 43036 29876 43092
rect 29708 43026 29764 43036
rect 29596 42980 29652 42990
rect 29596 42886 29652 42924
rect 29820 42866 29876 43036
rect 29820 42814 29822 42866
rect 29874 42814 29876 42866
rect 29820 42802 29876 42814
rect 29820 41972 29876 41982
rect 29820 41878 29876 41916
rect 29596 41746 29652 41758
rect 29596 41694 29598 41746
rect 29650 41694 29652 41746
rect 29596 41188 29652 41694
rect 29596 41186 29764 41188
rect 29596 41134 29598 41186
rect 29650 41134 29764 41186
rect 29596 41132 29764 41134
rect 29596 41122 29652 41132
rect 29708 40628 29764 41132
rect 29708 40534 29764 40572
rect 29372 39842 29540 39844
rect 29372 39790 29374 39842
rect 29426 39790 29540 39842
rect 29372 39788 29540 39790
rect 29596 40516 29652 40526
rect 29596 39842 29652 40460
rect 29596 39790 29598 39842
rect 29650 39790 29652 39842
rect 29372 39778 29428 39788
rect 29596 39778 29652 39790
rect 29820 40292 29876 40302
rect 29148 39620 29204 39630
rect 29148 39526 29204 39564
rect 29708 39506 29764 39518
rect 29708 39454 29710 39506
rect 29762 39454 29764 39506
rect 29260 39396 29316 39406
rect 29260 38834 29316 39340
rect 29260 38782 29262 38834
rect 29314 38782 29316 38834
rect 29260 38770 29316 38782
rect 29484 38836 29540 38874
rect 29708 38836 29764 39454
rect 29484 38770 29540 38780
rect 29596 38780 29764 38836
rect 29596 38668 29652 38780
rect 29260 38612 29316 38622
rect 29036 38434 29092 38444
rect 29148 38556 29260 38612
rect 28588 38052 28644 38062
rect 29036 38052 29092 38062
rect 28588 37958 28644 37996
rect 28924 38050 29092 38052
rect 28924 37998 29038 38050
rect 29090 37998 29092 38050
rect 28924 37996 29092 37998
rect 28924 37828 28980 37996
rect 29036 37986 29092 37996
rect 28924 37762 28980 37772
rect 28476 37266 28532 37436
rect 28476 37214 28478 37266
rect 28530 37214 28532 37266
rect 28476 37202 28532 37214
rect 28588 37380 28644 37390
rect 28588 37044 28644 37324
rect 28924 37268 28980 37278
rect 28924 37174 28980 37212
rect 29148 37156 29204 38556
rect 29260 38546 29316 38556
rect 29372 38612 29652 38668
rect 29260 38052 29316 38062
rect 29260 37958 29316 37996
rect 29372 38050 29428 38612
rect 29372 37998 29374 38050
rect 29426 37998 29428 38050
rect 29260 37380 29316 37390
rect 29372 37380 29428 37998
rect 29316 37324 29428 37380
rect 29484 38052 29540 38062
rect 29260 37314 29316 37324
rect 29148 37154 29428 37156
rect 29148 37102 29150 37154
rect 29202 37102 29428 37154
rect 29148 37100 29428 37102
rect 29148 37090 29204 37100
rect 28140 36764 28420 36820
rect 28476 36988 28644 37044
rect 28140 36596 28196 36764
rect 28140 36540 28308 36596
rect 28252 36482 28308 36540
rect 28252 36430 28254 36482
rect 28306 36430 28308 36482
rect 28140 36372 28196 36382
rect 28140 36278 28196 36316
rect 28252 36036 28308 36430
rect 28252 35970 28308 35980
rect 28364 35924 28420 35934
rect 28364 35830 28420 35868
rect 28140 33572 28196 33582
rect 28028 33516 28140 33572
rect 28140 33506 28196 33516
rect 27580 33406 27582 33458
rect 27634 33406 27636 33458
rect 27580 33394 27636 33406
rect 26684 33348 26740 33358
rect 26572 33346 26740 33348
rect 26572 33294 26686 33346
rect 26738 33294 26740 33346
rect 26572 33292 26740 33294
rect 26684 33282 26740 33292
rect 27020 33236 27076 33246
rect 27020 33142 27076 33180
rect 26908 33122 26964 33134
rect 26908 33070 26910 33122
rect 26962 33070 26964 33122
rect 26908 32676 26964 33070
rect 26908 32610 26964 32620
rect 26684 32564 26740 32574
rect 26348 32562 26740 32564
rect 26348 32510 26686 32562
rect 26738 32510 26740 32562
rect 26348 32508 26740 32510
rect 26684 32498 26740 32508
rect 26124 31714 26180 31724
rect 28476 31780 28532 36988
rect 29260 36932 29316 36942
rect 29148 36820 29204 36830
rect 29148 36482 29204 36764
rect 29260 36594 29316 36876
rect 29260 36542 29262 36594
rect 29314 36542 29316 36594
rect 29260 36530 29316 36542
rect 29148 36430 29150 36482
rect 29202 36430 29204 36482
rect 28812 36036 28868 36046
rect 28812 35922 28868 35980
rect 28812 35870 28814 35922
rect 28866 35870 28868 35922
rect 28812 35308 28868 35870
rect 28700 35252 28868 35308
rect 29148 35308 29204 36430
rect 29372 35924 29428 37100
rect 29484 36706 29540 37996
rect 29708 37940 29764 37950
rect 29708 37846 29764 37884
rect 29708 37380 29764 37390
rect 29820 37380 29876 40236
rect 29932 39620 29988 43484
rect 30156 42756 30212 42766
rect 30044 42642 30100 42654
rect 30044 42590 30046 42642
rect 30098 42590 30100 42642
rect 30044 41412 30100 42590
rect 30156 42530 30212 42700
rect 30156 42478 30158 42530
rect 30210 42478 30212 42530
rect 30156 42466 30212 42478
rect 30268 42194 30324 46284
rect 30380 45890 30436 45902
rect 30380 45838 30382 45890
rect 30434 45838 30436 45890
rect 30380 45780 30436 45838
rect 30380 45714 30436 45724
rect 30492 45780 30548 45790
rect 30492 45778 30660 45780
rect 30492 45726 30494 45778
rect 30546 45726 30660 45778
rect 30492 45724 30660 45726
rect 30492 45714 30548 45724
rect 30492 45444 30548 45454
rect 30380 43540 30436 43550
rect 30380 43446 30436 43484
rect 30380 42756 30436 42766
rect 30380 42662 30436 42700
rect 30268 42142 30270 42194
rect 30322 42142 30324 42194
rect 30268 41746 30324 42142
rect 30492 42196 30548 45388
rect 30604 45218 30660 45724
rect 30604 45166 30606 45218
rect 30658 45166 30660 45218
rect 30604 45154 30660 45166
rect 30716 45106 30772 48524
rect 30828 46340 30884 48748
rect 30828 46274 30884 46284
rect 30716 45054 30718 45106
rect 30770 45054 30772 45106
rect 30604 44324 30660 44334
rect 30604 44230 30660 44268
rect 30716 43764 30772 45054
rect 30940 44548 30996 49420
rect 31052 48356 31108 49532
rect 31164 49364 31220 49374
rect 31164 48356 31220 49308
rect 31276 48804 31332 48814
rect 31500 48804 31556 48814
rect 31276 48802 31556 48804
rect 31276 48750 31278 48802
rect 31330 48750 31502 48802
rect 31554 48750 31556 48802
rect 31276 48748 31556 48750
rect 31276 48738 31332 48748
rect 31500 48580 31556 48748
rect 31612 48804 31668 48814
rect 31612 48710 31668 48748
rect 31724 48804 31780 48814
rect 31836 48804 31892 49758
rect 31948 49028 32004 49038
rect 31948 48914 32004 48972
rect 31948 48862 31950 48914
rect 32002 48862 32004 48914
rect 31948 48850 32004 48862
rect 31724 48802 31892 48804
rect 31724 48750 31726 48802
rect 31778 48750 31892 48802
rect 31724 48748 31892 48750
rect 31724 48738 31780 48748
rect 31500 48524 31668 48580
rect 31500 48356 31556 48366
rect 31164 48354 31556 48356
rect 31164 48302 31502 48354
rect 31554 48302 31556 48354
rect 31164 48300 31556 48302
rect 31052 48290 31108 48300
rect 31500 48290 31556 48300
rect 31052 48132 31108 48142
rect 31052 48038 31108 48076
rect 31164 47684 31220 47694
rect 31164 47458 31220 47628
rect 31388 47572 31444 47582
rect 31388 47478 31444 47516
rect 31164 47406 31166 47458
rect 31218 47406 31220 47458
rect 31164 47394 31220 47406
rect 31388 46676 31444 46686
rect 31276 45890 31332 45902
rect 31276 45838 31278 45890
rect 31330 45838 31332 45890
rect 31276 45330 31332 45838
rect 31388 45668 31444 46620
rect 31500 45892 31556 45902
rect 31500 45798 31556 45836
rect 31388 45612 31556 45668
rect 31276 45278 31278 45330
rect 31330 45278 31332 45330
rect 31276 45266 31332 45278
rect 31388 45218 31444 45230
rect 31388 45166 31390 45218
rect 31442 45166 31444 45218
rect 31164 45108 31220 45118
rect 31164 45014 31220 45052
rect 30828 44492 30996 44548
rect 31388 44548 31444 45166
rect 30828 43876 30884 44492
rect 31388 44482 31444 44492
rect 31164 44436 31220 44446
rect 30940 44324 30996 44334
rect 30940 44098 30996 44268
rect 30940 44046 30942 44098
rect 30994 44046 30996 44098
rect 30940 44034 30996 44046
rect 31052 44210 31108 44222
rect 31052 44158 31054 44210
rect 31106 44158 31108 44210
rect 30828 43820 30996 43876
rect 30716 43708 30884 43764
rect 30604 43652 30660 43662
rect 30604 42756 30660 43596
rect 30828 43650 30884 43708
rect 30828 43598 30830 43650
rect 30882 43598 30884 43650
rect 30716 43540 30772 43550
rect 30716 42978 30772 43484
rect 30716 42926 30718 42978
rect 30770 42926 30772 42978
rect 30716 42914 30772 42926
rect 30828 42980 30884 43598
rect 30828 42914 30884 42924
rect 30604 42700 30884 42756
rect 30604 42530 30660 42542
rect 30604 42478 30606 42530
rect 30658 42478 30660 42530
rect 30604 42420 30660 42478
rect 30604 42354 30660 42364
rect 30492 42140 30772 42196
rect 30492 41972 30548 41982
rect 30268 41694 30270 41746
rect 30322 41694 30324 41746
rect 30268 41682 30324 41694
rect 30380 41970 30548 41972
rect 30380 41918 30494 41970
rect 30546 41918 30548 41970
rect 30380 41916 30548 41918
rect 30044 41298 30100 41356
rect 30044 41246 30046 41298
rect 30098 41246 30100 41298
rect 30044 41234 30100 41246
rect 30380 40964 30436 41916
rect 30492 41906 30548 41916
rect 30604 41972 30660 41982
rect 30604 41186 30660 41916
rect 30604 41134 30606 41186
rect 30658 41134 30660 41186
rect 30604 41122 30660 41134
rect 30268 40908 30436 40964
rect 30268 40852 30324 40908
rect 30156 40796 30324 40852
rect 30156 40292 30212 40796
rect 30268 40628 30324 40638
rect 30604 40628 30660 40638
rect 30716 40628 30772 42140
rect 30828 42194 30884 42700
rect 30828 42142 30830 42194
rect 30882 42142 30884 42194
rect 30828 42130 30884 42142
rect 30828 41972 30884 41982
rect 30828 41074 30884 41916
rect 30828 41022 30830 41074
rect 30882 41022 30884 41074
rect 30828 41010 30884 41022
rect 30268 40626 30772 40628
rect 30268 40574 30270 40626
rect 30322 40574 30606 40626
rect 30658 40574 30772 40626
rect 30268 40572 30772 40574
rect 30828 40628 30884 40638
rect 30268 40562 30324 40572
rect 30604 40562 30660 40572
rect 30828 40534 30884 40572
rect 30156 40226 30212 40236
rect 30492 40402 30548 40414
rect 30492 40350 30494 40402
rect 30546 40350 30548 40402
rect 29932 39554 29988 39564
rect 30492 38668 30548 40350
rect 30492 38612 30884 38668
rect 30156 38164 30212 38174
rect 30156 38070 30212 38108
rect 30156 37716 30212 37726
rect 29708 37378 29876 37380
rect 29708 37326 29710 37378
rect 29762 37326 29876 37378
rect 29708 37324 29876 37326
rect 30044 37660 30156 37716
rect 29708 37314 29764 37324
rect 29484 36654 29486 36706
rect 29538 36654 29540 36706
rect 29484 36036 29540 36654
rect 29484 35970 29540 35980
rect 29596 37268 29652 37278
rect 29596 35924 29652 37212
rect 30044 37266 30100 37660
rect 30156 37650 30212 37660
rect 30716 37492 30772 37502
rect 30716 37378 30772 37436
rect 30716 37326 30718 37378
rect 30770 37326 30772 37378
rect 30716 37314 30772 37326
rect 30044 37214 30046 37266
rect 30098 37214 30100 37266
rect 29932 36260 29988 36270
rect 29932 36166 29988 36204
rect 30044 36148 30100 37214
rect 30828 37268 30884 38612
rect 30940 38388 30996 43820
rect 31052 43764 31108 44158
rect 31052 43698 31108 43708
rect 31164 43540 31220 44380
rect 31052 43484 31220 43540
rect 31276 44210 31332 44222
rect 31276 44158 31278 44210
rect 31330 44158 31332 44210
rect 31052 42082 31108 43484
rect 31276 42644 31332 44158
rect 31388 43764 31444 43774
rect 31388 43650 31444 43708
rect 31388 43598 31390 43650
rect 31442 43598 31444 43650
rect 31388 43586 31444 43598
rect 31276 42578 31332 42588
rect 31500 42642 31556 45612
rect 31612 43988 31668 48524
rect 31724 47684 31780 47694
rect 31724 47590 31780 47628
rect 31724 47348 31780 47358
rect 31836 47348 31892 48748
rect 31948 48356 32004 48366
rect 31948 47458 32004 48300
rect 31948 47406 31950 47458
rect 32002 47406 32004 47458
rect 31948 47394 32004 47406
rect 32060 48132 32116 48142
rect 31780 47292 31892 47348
rect 31724 47282 31780 47292
rect 32060 47236 32116 48076
rect 31724 46562 31780 46574
rect 31724 46510 31726 46562
rect 31778 46510 31780 46562
rect 31724 45556 31780 46510
rect 31724 45490 31780 45500
rect 31836 44324 31892 44334
rect 31836 44230 31892 44268
rect 31612 43922 31668 43932
rect 32060 43204 32116 47180
rect 32172 47012 32228 50428
rect 32508 50148 32564 50428
rect 32732 50418 32788 50428
rect 32844 50482 32900 50494
rect 32844 50430 32846 50482
rect 32898 50430 32900 50482
rect 32620 50372 32676 50382
rect 32620 50278 32676 50316
rect 32844 50372 32900 50430
rect 32844 50306 32900 50316
rect 32508 50082 32564 50092
rect 32396 49924 32452 49934
rect 32396 49830 32452 49868
rect 32508 49140 32564 49150
rect 32956 49140 33012 49150
rect 32508 49138 33012 49140
rect 32508 49086 32510 49138
rect 32562 49086 32958 49138
rect 33010 49086 33012 49138
rect 32508 49084 33012 49086
rect 32508 49074 32564 49084
rect 32956 49074 33012 49084
rect 32396 48804 32452 48814
rect 32620 48804 32676 48814
rect 32396 48710 32452 48748
rect 32508 48802 32676 48804
rect 32508 48750 32622 48802
rect 32674 48750 32676 48802
rect 32508 48748 32676 48750
rect 32508 47572 32564 48748
rect 32620 48738 32676 48748
rect 32844 48802 32900 48814
rect 32844 48750 32846 48802
rect 32898 48750 32900 48802
rect 32620 48130 32676 48142
rect 32620 48078 32622 48130
rect 32674 48078 32676 48130
rect 32620 47796 32676 48078
rect 32844 48132 32900 48750
rect 33068 48466 33124 52668
rect 33404 52164 33460 53228
rect 33516 52722 33572 55020
rect 33628 54740 33684 54750
rect 33628 54626 33684 54684
rect 33628 54574 33630 54626
rect 33682 54574 33684 54626
rect 33628 54180 33684 54574
rect 33628 54114 33684 54124
rect 33852 53730 33908 55246
rect 34300 55076 34356 55916
rect 34412 55524 34468 56252
rect 35308 55972 35364 55982
rect 35308 55878 35364 55916
rect 36092 55972 36148 55982
rect 36092 55878 36148 55916
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 34412 55468 35028 55524
rect 34412 55298 34468 55468
rect 34412 55246 34414 55298
rect 34466 55246 34468 55298
rect 34412 55234 34468 55246
rect 34860 55188 34916 55198
rect 34860 55094 34916 55132
rect 34300 55010 34356 55020
rect 34748 54740 34804 54750
rect 34524 54516 34580 54526
rect 34076 54514 34580 54516
rect 34076 54462 34526 54514
rect 34578 54462 34580 54514
rect 34076 54460 34580 54462
rect 33852 53678 33854 53730
rect 33906 53678 33908 53730
rect 33852 53508 33908 53678
rect 33628 53172 33684 53182
rect 33628 53078 33684 53116
rect 33516 52670 33518 52722
rect 33570 52670 33572 52722
rect 33516 52658 33572 52670
rect 33852 52722 33908 53452
rect 33964 54404 34020 54414
rect 33964 53172 34020 54348
rect 34076 53956 34132 54460
rect 34524 54450 34580 54460
rect 34076 53862 34132 53900
rect 34300 54180 34356 54190
rect 34300 53954 34356 54124
rect 34300 53902 34302 53954
rect 34354 53902 34356 53954
rect 34300 53890 34356 53902
rect 34748 53954 34804 54684
rect 34748 53902 34750 53954
rect 34802 53902 34804 53954
rect 34748 53890 34804 53902
rect 34860 54516 34916 54526
rect 34972 54516 35028 55468
rect 35980 55412 36036 55422
rect 35980 55298 36036 55356
rect 35980 55246 35982 55298
rect 36034 55246 36036 55298
rect 35980 55234 36036 55246
rect 36204 55298 36260 55310
rect 36204 55246 36206 55298
rect 36258 55246 36260 55298
rect 34860 54514 35028 54516
rect 34860 54462 34862 54514
rect 34914 54462 35028 54514
rect 34860 54460 35028 54462
rect 36092 54514 36148 54526
rect 36092 54462 36094 54514
rect 36146 54462 36148 54514
rect 34524 53620 34580 53630
rect 34076 53172 34132 53182
rect 33964 53170 34132 53172
rect 33964 53118 34078 53170
rect 34130 53118 34132 53170
rect 33964 53116 34132 53118
rect 34076 53106 34132 53116
rect 33852 52670 33854 52722
rect 33906 52670 33908 52722
rect 33852 52658 33908 52670
rect 34524 52834 34580 53564
rect 34860 53172 34916 54460
rect 35420 54404 35476 54414
rect 35420 54402 35588 54404
rect 35420 54350 35422 54402
rect 35474 54350 35588 54402
rect 35420 54348 35588 54350
rect 35420 54338 35476 54348
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 35420 53956 35476 53966
rect 35196 53844 35252 53854
rect 35196 53750 35252 53788
rect 35420 53842 35476 53900
rect 35420 53790 35422 53842
rect 35474 53790 35476 53842
rect 35420 53778 35476 53790
rect 35532 53730 35588 54348
rect 35532 53678 35534 53730
rect 35586 53678 35588 53730
rect 34860 53106 34916 53116
rect 35420 53172 35476 53182
rect 35420 53078 35476 53116
rect 34972 53060 35028 53070
rect 34972 52966 35028 53004
rect 34524 52782 34526 52834
rect 34578 52782 34580 52834
rect 34524 52724 34580 52782
rect 34524 52658 34580 52668
rect 34636 52722 34692 52734
rect 34636 52670 34638 52722
rect 34690 52670 34692 52722
rect 33852 52274 33908 52286
rect 33852 52222 33854 52274
rect 33906 52222 33908 52274
rect 33852 52164 33908 52222
rect 34300 52164 34356 52174
rect 33404 52162 33572 52164
rect 33404 52110 33406 52162
rect 33458 52110 33572 52162
rect 33404 52108 33572 52110
rect 33404 52098 33460 52108
rect 33180 51266 33236 51278
rect 33180 51214 33182 51266
rect 33234 51214 33236 51266
rect 33180 51044 33236 51214
rect 33180 50978 33236 50988
rect 33292 51156 33348 51166
rect 33292 50706 33348 51100
rect 33292 50654 33294 50706
rect 33346 50654 33348 50706
rect 33292 50642 33348 50654
rect 33516 50596 33572 52108
rect 33852 52162 34356 52164
rect 33852 52110 34302 52162
rect 34354 52110 34356 52162
rect 33852 52108 34356 52110
rect 33740 51604 33796 51614
rect 33740 51378 33796 51548
rect 33740 51326 33742 51378
rect 33794 51326 33796 51378
rect 33740 51314 33796 51326
rect 33740 50596 33796 50634
rect 33516 50540 33684 50596
rect 33516 50372 33572 50540
rect 33516 50306 33572 50316
rect 33628 50034 33684 50540
rect 33740 50530 33796 50540
rect 33852 50428 33908 52108
rect 34300 52098 34356 52108
rect 34524 52162 34580 52174
rect 34524 52110 34526 52162
rect 34578 52110 34580 52162
rect 34188 51378 34244 51390
rect 34188 51326 34190 51378
rect 34242 51326 34244 51378
rect 34188 50932 34244 51326
rect 34188 50596 34244 50876
rect 34188 50530 34244 50540
rect 34524 51266 34580 52110
rect 34524 51214 34526 51266
rect 34578 51214 34580 51266
rect 34524 50428 34580 51214
rect 33628 49982 33630 50034
rect 33682 49982 33684 50034
rect 33628 49970 33684 49982
rect 33740 50372 33908 50428
rect 34076 50372 34580 50428
rect 33516 49810 33572 49822
rect 33516 49758 33518 49810
rect 33570 49758 33572 49810
rect 33516 49250 33572 49758
rect 33516 49198 33518 49250
rect 33570 49198 33572 49250
rect 33516 49186 33572 49198
rect 33404 49028 33460 49038
rect 33404 48934 33460 48972
rect 33068 48414 33070 48466
rect 33122 48414 33124 48466
rect 33068 48402 33124 48414
rect 33628 48354 33684 48366
rect 33628 48302 33630 48354
rect 33682 48302 33684 48354
rect 32844 48066 32900 48076
rect 32956 48244 33012 48254
rect 32844 47796 32900 47806
rect 32620 47740 32844 47796
rect 32172 46946 32228 46956
rect 32284 47516 32564 47572
rect 32844 47570 32900 47740
rect 32844 47518 32846 47570
rect 32898 47518 32900 47570
rect 32284 46340 32340 47516
rect 32844 47506 32900 47518
rect 32060 43138 32116 43148
rect 32172 46284 32340 46340
rect 32396 47348 32452 47358
rect 32060 42980 32116 42990
rect 31836 42756 31892 42766
rect 31836 42662 31892 42700
rect 31500 42590 31502 42642
rect 31554 42590 31556 42642
rect 31164 42532 31220 42542
rect 31164 42438 31220 42476
rect 31052 42030 31054 42082
rect 31106 42030 31108 42082
rect 31052 40404 31108 42030
rect 31164 42084 31220 42094
rect 31164 41970 31220 42028
rect 31164 41918 31166 41970
rect 31218 41918 31220 41970
rect 31164 41906 31220 41918
rect 31500 41972 31556 42590
rect 31612 42532 31668 42542
rect 31612 42438 31668 42476
rect 31500 41906 31556 41916
rect 31276 41412 31332 41422
rect 31164 41356 31276 41412
rect 31164 41074 31220 41356
rect 31276 41346 31332 41356
rect 31388 41300 31444 41310
rect 31388 41188 31444 41244
rect 31164 41022 31166 41074
rect 31218 41022 31220 41074
rect 31164 41010 31220 41022
rect 31276 41132 31444 41188
rect 31500 41188 31556 41226
rect 31276 40514 31332 41132
rect 31500 41122 31556 41132
rect 31500 40964 31556 40974
rect 31276 40462 31278 40514
rect 31330 40462 31332 40514
rect 31276 40450 31332 40462
rect 31388 40962 31556 40964
rect 31388 40910 31502 40962
rect 31554 40910 31556 40962
rect 31388 40908 31556 40910
rect 31164 40404 31220 40414
rect 31052 40402 31220 40404
rect 31052 40350 31166 40402
rect 31218 40350 31220 40402
rect 31052 40348 31220 40350
rect 31164 40292 31220 40348
rect 31164 40236 31332 40292
rect 30940 38322 30996 38332
rect 31164 38052 31220 38062
rect 31164 37958 31220 37996
rect 30940 37268 30996 37278
rect 30828 37266 30996 37268
rect 30828 37214 30942 37266
rect 30994 37214 30996 37266
rect 30828 37212 30996 37214
rect 30156 37154 30212 37166
rect 30156 37102 30158 37154
rect 30210 37102 30212 37154
rect 30156 37044 30212 37102
rect 30156 36978 30212 36988
rect 30380 36708 30436 36718
rect 30380 36594 30436 36652
rect 30380 36542 30382 36594
rect 30434 36542 30436 36594
rect 30380 36530 30436 36542
rect 30716 36372 30772 36382
rect 30716 36278 30772 36316
rect 30044 36092 30324 36148
rect 29708 35924 29764 35934
rect 29596 35922 29764 35924
rect 29596 35870 29710 35922
rect 29762 35870 29764 35922
rect 29596 35868 29764 35870
rect 29372 35858 29428 35868
rect 29708 35858 29764 35868
rect 30156 35922 30212 35934
rect 30156 35870 30158 35922
rect 30210 35870 30212 35922
rect 29484 35810 29540 35822
rect 29484 35758 29486 35810
rect 29538 35758 29540 35810
rect 29372 35700 29428 35710
rect 29372 35606 29428 35644
rect 29148 35252 29316 35308
rect 28700 35026 28756 35252
rect 28700 34974 28702 35026
rect 28754 34974 28756 35026
rect 28700 34916 28756 34974
rect 28700 34850 28756 34860
rect 29148 35140 29204 35150
rect 29148 34916 29204 35084
rect 29260 35028 29316 35252
rect 29484 35252 29540 35758
rect 29484 35186 29540 35196
rect 29708 35700 29764 35710
rect 29820 35700 29876 35710
rect 29764 35698 29876 35700
rect 29764 35646 29822 35698
rect 29874 35646 29876 35698
rect 29764 35644 29876 35646
rect 29260 34972 29540 35028
rect 29148 34914 29316 34916
rect 29148 34862 29150 34914
rect 29202 34862 29316 34914
rect 29148 34860 29316 34862
rect 29148 34850 29204 34860
rect 29260 34242 29316 34860
rect 29484 34802 29540 34972
rect 29484 34750 29486 34802
rect 29538 34750 29540 34802
rect 29484 34692 29540 34750
rect 29484 34626 29540 34636
rect 29260 34190 29262 34242
rect 29314 34190 29316 34242
rect 29260 34178 29316 34190
rect 29708 34130 29764 35644
rect 29820 35634 29876 35644
rect 29708 34078 29710 34130
rect 29762 34078 29764 34130
rect 29708 34066 29764 34078
rect 30044 35252 30100 35262
rect 30044 34130 30100 35196
rect 30156 34916 30212 35870
rect 30268 35810 30324 36092
rect 30268 35758 30270 35810
rect 30322 35758 30324 35810
rect 30268 35252 30324 35758
rect 30268 35186 30324 35196
rect 30380 35698 30436 35710
rect 30380 35646 30382 35698
rect 30434 35646 30436 35698
rect 30268 34916 30324 34926
rect 30156 34914 30324 34916
rect 30156 34862 30270 34914
rect 30322 34862 30324 34914
rect 30156 34860 30324 34862
rect 30268 34850 30324 34860
rect 30156 34580 30212 34590
rect 30156 34354 30212 34524
rect 30156 34302 30158 34354
rect 30210 34302 30212 34354
rect 30156 34290 30212 34302
rect 30380 34356 30436 35646
rect 30380 34290 30436 34300
rect 30492 34914 30548 34926
rect 30492 34862 30494 34914
rect 30546 34862 30548 34914
rect 30492 34244 30548 34862
rect 30604 34692 30660 34702
rect 30604 34354 30660 34636
rect 30604 34302 30606 34354
rect 30658 34302 30660 34354
rect 30604 34290 30660 34302
rect 30492 34178 30548 34188
rect 30044 34078 30046 34130
rect 30098 34078 30100 34130
rect 30044 34066 30100 34078
rect 30828 34020 30884 37212
rect 30940 37202 30996 37212
rect 31276 37156 31332 40236
rect 31388 38948 31444 40908
rect 31500 40898 31556 40908
rect 32060 40626 32116 42924
rect 32172 40852 32228 46284
rect 32284 46116 32340 46126
rect 32284 45890 32340 46060
rect 32284 45838 32286 45890
rect 32338 45838 32340 45890
rect 32284 45826 32340 45838
rect 32396 45890 32452 47292
rect 32956 46900 33012 48188
rect 32396 45838 32398 45890
rect 32450 45838 32452 45890
rect 32396 45826 32452 45838
rect 32508 46844 32956 46900
rect 32508 46674 32564 46844
rect 32956 46834 33012 46844
rect 33068 48242 33124 48254
rect 33068 48190 33070 48242
rect 33122 48190 33124 48242
rect 32508 46622 32510 46674
rect 32562 46622 32564 46674
rect 32508 45444 32564 46622
rect 32844 46116 32900 46126
rect 32844 46022 32900 46060
rect 33068 46004 33124 48190
rect 33516 48242 33572 48254
rect 33516 48190 33518 48242
rect 33570 48190 33572 48242
rect 33180 48130 33236 48142
rect 33180 48078 33182 48130
rect 33234 48078 33236 48130
rect 33180 47796 33236 48078
rect 33516 47796 33572 48190
rect 33180 47740 33348 47796
rect 33292 47460 33348 47740
rect 33404 47460 33460 47470
rect 33292 47458 33460 47460
rect 33292 47406 33406 47458
rect 33458 47406 33460 47458
rect 33292 47404 33460 47406
rect 33180 46900 33236 46910
rect 33180 46806 33236 46844
rect 32956 45948 33124 46004
rect 32732 45890 32788 45902
rect 32956 45892 33012 45948
rect 32732 45838 32734 45890
rect 32786 45838 32788 45890
rect 32508 45378 32564 45388
rect 32620 45668 32676 45678
rect 32508 45108 32564 45118
rect 32508 45014 32564 45052
rect 32284 44548 32340 44558
rect 32284 44322 32340 44492
rect 32620 44434 32676 45612
rect 32620 44382 32622 44434
rect 32674 44382 32676 44434
rect 32620 44370 32676 44382
rect 32732 44436 32788 45838
rect 32732 44370 32788 44380
rect 32844 45836 33012 45892
rect 32284 44270 32286 44322
rect 32338 44270 32340 44322
rect 32284 43876 32340 44270
rect 32284 43810 32340 43820
rect 32844 44322 32900 45836
rect 33068 45218 33124 45230
rect 33068 45166 33070 45218
rect 33122 45166 33124 45218
rect 33068 44436 33124 45166
rect 33068 44370 33124 44380
rect 32844 44270 32846 44322
rect 32898 44270 32900 44322
rect 32844 43764 32900 44270
rect 33068 44212 33124 44222
rect 33068 44118 33124 44156
rect 32844 43698 32900 43708
rect 33180 42980 33236 42990
rect 32396 42756 32452 42766
rect 32396 42662 32452 42700
rect 32508 42644 32564 42654
rect 32508 42550 32564 42588
rect 32732 42644 32788 42654
rect 32732 42550 32788 42588
rect 33180 42196 33236 42924
rect 32956 42194 33236 42196
rect 32956 42142 33182 42194
rect 33234 42142 33236 42194
rect 32956 42140 33236 42142
rect 32172 40786 32228 40796
rect 32620 41186 32676 41198
rect 32620 41134 32622 41186
rect 32674 41134 32676 41186
rect 32060 40574 32062 40626
rect 32114 40574 32116 40626
rect 31836 40516 31892 40526
rect 31724 40514 31892 40516
rect 31724 40462 31838 40514
rect 31890 40462 31892 40514
rect 31724 40460 31892 40462
rect 31500 40404 31556 40414
rect 31500 40310 31556 40348
rect 31724 40402 31780 40460
rect 31836 40450 31892 40460
rect 31724 40350 31726 40402
rect 31778 40350 31780 40402
rect 31724 40338 31780 40350
rect 31948 40404 32004 40414
rect 31724 40180 31780 40190
rect 31724 39730 31780 40124
rect 31948 39844 32004 40348
rect 32060 40180 32116 40574
rect 32172 40404 32228 40414
rect 32172 40402 32340 40404
rect 32172 40350 32174 40402
rect 32226 40350 32340 40402
rect 32172 40348 32340 40350
rect 32172 40338 32228 40348
rect 32060 40114 32116 40124
rect 31948 39788 32228 39844
rect 31724 39678 31726 39730
rect 31778 39678 31780 39730
rect 31724 39666 31780 39678
rect 31948 39620 32004 39630
rect 31724 39284 31780 39294
rect 31388 38892 31668 38948
rect 31612 38668 31668 38892
rect 31724 38834 31780 39228
rect 31724 38782 31726 38834
rect 31778 38782 31780 38834
rect 31724 38770 31780 38782
rect 31948 38834 32004 39564
rect 32060 39618 32116 39630
rect 32060 39566 32062 39618
rect 32114 39566 32116 39618
rect 32060 39172 32116 39566
rect 32060 39106 32116 39116
rect 31948 38782 31950 38834
rect 32002 38782 32004 38834
rect 31948 38770 32004 38782
rect 32060 38724 32116 38734
rect 31612 38612 31780 38668
rect 31724 38050 31780 38612
rect 31724 37998 31726 38050
rect 31778 37998 31780 38050
rect 31724 37986 31780 37998
rect 32060 38050 32116 38668
rect 32172 38162 32228 39788
rect 32284 39732 32340 40348
rect 32284 39506 32340 39676
rect 32284 39454 32286 39506
rect 32338 39454 32340 39506
rect 32284 39442 32340 39454
rect 32172 38110 32174 38162
rect 32226 38110 32228 38162
rect 32172 38098 32228 38110
rect 32284 38834 32340 38846
rect 32284 38782 32286 38834
rect 32338 38782 32340 38834
rect 32060 37998 32062 38050
rect 32114 37998 32116 38050
rect 32060 37986 32116 37998
rect 32284 37604 32340 38782
rect 32508 38724 32564 38762
rect 32060 37548 32340 37604
rect 32396 38610 32452 38622
rect 32396 38558 32398 38610
rect 32450 38558 32452 38610
rect 31276 37090 31332 37100
rect 31948 37268 32004 37278
rect 31948 37154 32004 37212
rect 31948 37102 31950 37154
rect 32002 37102 32004 37154
rect 31948 37090 32004 37102
rect 32060 37266 32116 37548
rect 32172 37380 32228 37390
rect 32172 37286 32228 37324
rect 32060 37214 32062 37266
rect 32114 37214 32116 37266
rect 32060 36932 32116 37214
rect 32284 37268 32340 37278
rect 32396 37268 32452 38558
rect 32508 37492 32564 38668
rect 32620 37716 32676 41134
rect 32844 38500 32900 38510
rect 32844 38050 32900 38444
rect 32844 37998 32846 38050
rect 32898 37998 32900 38050
rect 32844 37986 32900 37998
rect 32620 37650 32676 37660
rect 32508 37436 32676 37492
rect 32396 37212 32564 37268
rect 31052 36596 31108 36606
rect 31500 36596 31556 36606
rect 31052 36594 31444 36596
rect 31052 36542 31054 36594
rect 31106 36542 31444 36594
rect 31052 36540 31444 36542
rect 31052 36530 31108 36540
rect 31388 36482 31444 36540
rect 31388 36430 31390 36482
rect 31442 36430 31444 36482
rect 31388 36418 31444 36430
rect 30940 36372 30996 36382
rect 30940 36278 30996 36316
rect 31052 35252 31108 35262
rect 30940 35026 30996 35038
rect 30940 34974 30942 35026
rect 30994 34974 30996 35026
rect 30940 34916 30996 34974
rect 30940 34850 30996 34860
rect 31052 34914 31108 35196
rect 31276 35140 31332 35150
rect 31500 35140 31556 36540
rect 32060 36372 32116 36876
rect 32060 36306 32116 36316
rect 32172 37156 32228 37166
rect 31276 35138 31556 35140
rect 31276 35086 31278 35138
rect 31330 35086 31556 35138
rect 31276 35084 31556 35086
rect 31276 35074 31332 35084
rect 31052 34862 31054 34914
rect 31106 34862 31108 34914
rect 30380 33964 30884 34020
rect 31052 34018 31108 34862
rect 32060 35028 32116 35038
rect 32060 34690 32116 34972
rect 32172 34916 32228 37100
rect 32284 35140 32340 37212
rect 32396 37044 32452 37054
rect 32396 36482 32452 36988
rect 32396 36430 32398 36482
rect 32450 36430 32452 36482
rect 32396 36418 32452 36430
rect 32508 36148 32564 37212
rect 32620 36370 32676 37436
rect 32956 36708 33012 42140
rect 33180 42130 33236 42140
rect 33292 38668 33348 47404
rect 33404 47394 33460 47404
rect 33516 47236 33572 47740
rect 33628 47460 33684 48302
rect 33740 47572 33796 50372
rect 33852 49810 33908 49822
rect 33852 49758 33854 49810
rect 33906 49758 33908 49810
rect 33852 49588 33908 49758
rect 33964 49588 34020 49598
rect 33852 49586 34020 49588
rect 33852 49534 33966 49586
rect 34018 49534 34020 49586
rect 33852 49532 34020 49534
rect 33964 49522 34020 49532
rect 33740 47506 33796 47516
rect 33628 47366 33684 47404
rect 33740 47346 33796 47358
rect 33740 47294 33742 47346
rect 33794 47294 33796 47346
rect 33740 47236 33796 47294
rect 33516 47180 34020 47236
rect 33628 47012 33684 47022
rect 33404 45220 33460 45230
rect 33404 45126 33460 45164
rect 33404 44772 33460 44782
rect 33404 44100 33460 44716
rect 33404 43762 33460 44044
rect 33404 43710 33406 43762
rect 33458 43710 33460 43762
rect 33404 43652 33460 43710
rect 33404 43586 33460 43596
rect 33628 44100 33684 46956
rect 33852 46564 33908 46574
rect 33852 46114 33908 46508
rect 33852 46062 33854 46114
rect 33906 46062 33908 46114
rect 33852 46004 33908 46062
rect 33404 43204 33460 43214
rect 33404 39508 33460 43148
rect 33628 42196 33684 44044
rect 33740 46002 33908 46004
rect 33740 45950 33854 46002
rect 33906 45950 33908 46002
rect 33740 45948 33908 45950
rect 33740 43762 33796 45948
rect 33852 45938 33908 45948
rect 33740 43710 33742 43762
rect 33794 43710 33796 43762
rect 33740 43428 33796 43710
rect 33740 43362 33796 43372
rect 33852 45108 33908 45118
rect 33852 44210 33908 45052
rect 33964 44548 34020 47180
rect 34076 46228 34132 50372
rect 34300 49810 34356 49822
rect 34300 49758 34302 49810
rect 34354 49758 34356 49810
rect 34300 49698 34356 49758
rect 34300 49646 34302 49698
rect 34354 49646 34356 49698
rect 34300 49634 34356 49646
rect 34636 49252 34692 52670
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 34860 52164 34916 52174
rect 34860 51938 34916 52108
rect 34860 51886 34862 51938
rect 34914 51886 34916 51938
rect 34860 51874 34916 51886
rect 35196 52162 35252 52174
rect 35196 52110 35198 52162
rect 35250 52110 35252 52162
rect 35196 51604 35252 52110
rect 35420 52164 35476 52174
rect 35420 52070 35476 52108
rect 35196 51538 35252 51548
rect 34860 51492 34916 51502
rect 34860 51398 34916 51436
rect 35308 51492 35364 51502
rect 35532 51492 35588 53678
rect 36092 53620 36148 54462
rect 36204 53844 36260 55246
rect 36204 53778 36260 53788
rect 35980 53508 36036 53518
rect 35980 53414 36036 53452
rect 35308 51490 35588 51492
rect 35308 51438 35310 51490
rect 35362 51438 35588 51490
rect 35308 51436 35588 51438
rect 35644 52388 35700 52398
rect 35308 51426 35364 51436
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 35196 50708 35252 50718
rect 35196 49922 35252 50652
rect 35644 50484 35700 52332
rect 35756 52388 35812 52398
rect 36092 52388 36148 53564
rect 36316 52724 36372 57708
rect 38556 57540 38612 57550
rect 37100 56756 37156 56766
rect 36988 56084 37044 56094
rect 36988 55990 37044 56028
rect 36540 55970 36596 55982
rect 36540 55918 36542 55970
rect 36594 55918 36596 55970
rect 36540 55524 36596 55918
rect 36540 55458 36596 55468
rect 36428 55188 36484 55198
rect 36428 55094 36484 55132
rect 36652 55076 36708 55086
rect 36652 54514 36708 55020
rect 36652 54462 36654 54514
rect 36706 54462 36708 54514
rect 36652 54450 36708 54462
rect 36988 54852 37044 54862
rect 36764 53844 36820 53854
rect 36428 53506 36484 53518
rect 36428 53454 36430 53506
rect 36482 53454 36484 53506
rect 36428 52948 36484 53454
rect 36428 52882 36484 52892
rect 36316 52668 36484 52724
rect 35756 52386 36148 52388
rect 35756 52334 35758 52386
rect 35810 52334 36148 52386
rect 35756 52332 36148 52334
rect 35756 52322 35812 52332
rect 36316 50594 36372 50606
rect 36316 50542 36318 50594
rect 36370 50542 36372 50594
rect 35756 50484 35812 50522
rect 35644 50482 35812 50484
rect 35644 50430 35758 50482
rect 35810 50430 35812 50482
rect 35644 50428 35812 50430
rect 36316 50484 36372 50542
rect 35196 49870 35198 49922
rect 35250 49870 35252 49922
rect 35196 49858 35252 49870
rect 35756 50372 36148 50428
rect 36316 50418 36372 50428
rect 35420 49812 35476 49822
rect 35420 49718 35476 49756
rect 34972 49700 35028 49710
rect 34972 49606 35028 49644
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 34300 49196 34692 49252
rect 34188 47348 34244 47358
rect 34188 47254 34244 47292
rect 34076 46162 34132 46172
rect 34300 45892 34356 49196
rect 34412 49028 34468 49038
rect 34412 48242 34468 48972
rect 34748 48802 34804 48814
rect 34748 48750 34750 48802
rect 34802 48750 34804 48802
rect 34412 48190 34414 48242
rect 34466 48190 34468 48242
rect 34412 48178 34468 48190
rect 34524 48466 34580 48478
rect 34524 48414 34526 48466
rect 34578 48414 34580 48466
rect 34524 48244 34580 48414
rect 34748 48468 34804 48750
rect 34748 48412 35140 48468
rect 35084 48354 35140 48412
rect 35084 48302 35086 48354
rect 35138 48302 35140 48354
rect 34972 48244 35028 48254
rect 34524 48242 35028 48244
rect 34524 48190 34974 48242
rect 35026 48190 35028 48242
rect 34524 48188 35028 48190
rect 34972 46786 35028 48188
rect 35084 47572 35140 48302
rect 35532 48130 35588 48142
rect 35532 48078 35534 48130
rect 35586 48078 35588 48130
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 35308 47572 35364 47582
rect 35084 47516 35252 47572
rect 35084 47346 35140 47358
rect 35084 47294 35086 47346
rect 35138 47294 35140 47346
rect 35084 46898 35140 47294
rect 35084 46846 35086 46898
rect 35138 46846 35140 46898
rect 35084 46834 35140 46846
rect 34972 46734 34974 46786
rect 35026 46734 35028 46786
rect 34972 46722 35028 46734
rect 35196 46674 35252 47516
rect 35196 46622 35198 46674
rect 35250 46622 35252 46674
rect 34636 46564 34692 46574
rect 35196 46564 35252 46622
rect 34636 46562 35252 46564
rect 34636 46510 34638 46562
rect 34690 46510 35252 46562
rect 34636 46508 35252 46510
rect 35308 47458 35364 47516
rect 35308 47406 35310 47458
rect 35362 47406 35364 47458
rect 34636 46498 34692 46508
rect 34300 45826 34356 45836
rect 34636 46114 34692 46126
rect 34636 46062 34638 46114
rect 34690 46062 34692 46114
rect 34300 45666 34356 45678
rect 34300 45614 34302 45666
rect 34354 45614 34356 45666
rect 34076 45220 34132 45230
rect 34076 45126 34132 45164
rect 34300 45106 34356 45614
rect 34300 45054 34302 45106
rect 34354 45054 34356 45106
rect 34300 44772 34356 45054
rect 34300 44706 34356 44716
rect 34412 45330 34468 45342
rect 34412 45278 34414 45330
rect 34466 45278 34468 45330
rect 33964 44492 34356 44548
rect 33852 44158 33854 44210
rect 33906 44158 33908 44210
rect 33740 42196 33796 42206
rect 33628 42140 33740 42196
rect 33740 42102 33796 42140
rect 33628 41746 33684 41758
rect 33628 41694 33630 41746
rect 33682 41694 33684 41746
rect 33628 41412 33684 41694
rect 33628 41186 33684 41356
rect 33628 41134 33630 41186
rect 33682 41134 33684 41186
rect 33628 41122 33684 41134
rect 33852 40068 33908 44158
rect 33964 44322 34020 44334
rect 33964 44270 33966 44322
rect 34018 44270 34020 44322
rect 33964 43764 34020 44270
rect 33964 43698 34020 43708
rect 34188 43988 34244 43998
rect 34188 41972 34244 43932
rect 34300 42980 34356 44492
rect 34412 43762 34468 45278
rect 34636 45218 34692 46062
rect 34636 45166 34638 45218
rect 34690 45166 34692 45218
rect 34636 45154 34692 45166
rect 34524 44996 34580 45006
rect 34524 44434 34580 44940
rect 34748 44884 34804 46508
rect 35308 46452 35364 47406
rect 35532 47012 35588 48078
rect 35756 48130 35812 50372
rect 36092 50034 36148 50372
rect 36092 49982 36094 50034
rect 36146 49982 36148 50034
rect 36092 49970 36148 49982
rect 36316 49812 36372 49822
rect 35980 48244 36036 48254
rect 35756 48078 35758 48130
rect 35810 48078 35812 48130
rect 35756 48066 35812 48078
rect 35868 48242 36036 48244
rect 35868 48190 35982 48242
rect 36034 48190 36036 48242
rect 35868 48188 36036 48190
rect 35756 47684 35812 47694
rect 35756 47590 35812 47628
rect 35532 46946 35588 46956
rect 35868 47348 35924 48188
rect 35980 48178 36036 48188
rect 35532 46788 35588 46798
rect 35868 46788 35924 47292
rect 35532 46786 35924 46788
rect 35532 46734 35534 46786
rect 35586 46734 35924 46786
rect 35532 46732 35924 46734
rect 35980 47684 36036 47694
rect 35532 46722 35588 46732
rect 35980 46674 36036 47628
rect 36092 47236 36148 47246
rect 36092 47234 36260 47236
rect 36092 47182 36094 47234
rect 36146 47182 36260 47234
rect 36092 47180 36260 47182
rect 36092 47170 36148 47180
rect 35980 46622 35982 46674
rect 36034 46622 36036 46674
rect 35980 46610 36036 46622
rect 36204 46676 36260 47180
rect 36204 46610 36260 46620
rect 36316 46786 36372 49756
rect 36428 49140 36484 52668
rect 36764 51380 36820 53788
rect 36876 53730 36932 53742
rect 36876 53678 36878 53730
rect 36930 53678 36932 53730
rect 36876 53620 36932 53678
rect 36876 53554 36932 53564
rect 36988 53172 37044 54796
rect 36988 53106 37044 53116
rect 36988 52836 37044 52846
rect 36876 51380 36932 51390
rect 36764 51378 36932 51380
rect 36764 51326 36878 51378
rect 36930 51326 36932 51378
rect 36764 51324 36932 51326
rect 36428 49046 36484 49084
rect 36540 51266 36596 51278
rect 36540 51214 36542 51266
rect 36594 51214 36596 51266
rect 36316 46734 36318 46786
rect 36370 46734 36372 46786
rect 36316 46452 36372 46734
rect 35084 46396 35364 46452
rect 35532 46396 36372 46452
rect 34748 44818 34804 44828
rect 34860 45778 34916 45790
rect 34860 45726 34862 45778
rect 34914 45726 34916 45778
rect 34524 44382 34526 44434
rect 34578 44382 34580 44434
rect 34524 44370 34580 44382
rect 34748 44436 34804 44446
rect 34524 44212 34580 44222
rect 34748 44212 34804 44380
rect 34524 44210 34804 44212
rect 34524 44158 34526 44210
rect 34578 44158 34804 44210
rect 34524 44156 34804 44158
rect 34524 44146 34580 44156
rect 34412 43710 34414 43762
rect 34466 43710 34468 43762
rect 34412 43698 34468 43710
rect 34524 43876 34580 43886
rect 34356 42924 34468 42980
rect 34300 42914 34356 42924
rect 34412 42866 34468 42924
rect 34412 42814 34414 42866
rect 34466 42814 34468 42866
rect 34412 42802 34468 42814
rect 34188 41878 34244 41916
rect 34300 42754 34356 42766
rect 34300 42702 34302 42754
rect 34354 42702 34356 42754
rect 34300 41746 34356 42702
rect 34300 41694 34302 41746
rect 34354 41694 34356 41746
rect 34300 41682 34356 41694
rect 34412 41524 34468 41534
rect 33852 40002 33908 40012
rect 34076 41298 34132 41310
rect 34076 41246 34078 41298
rect 34130 41246 34132 41298
rect 34076 41076 34132 41246
rect 34412 41188 34468 41468
rect 33516 39732 33572 39742
rect 33516 39638 33572 39676
rect 33404 39452 33908 39508
rect 33516 39172 33572 39182
rect 33404 39060 33460 39070
rect 33404 38966 33460 39004
rect 33516 38836 33572 39116
rect 33180 38612 33348 38668
rect 33404 38780 33572 38836
rect 33852 39058 33908 39452
rect 33852 39006 33854 39058
rect 33906 39006 33908 39058
rect 33068 38052 33124 38062
rect 33068 37958 33124 37996
rect 33068 37378 33124 37390
rect 33068 37326 33070 37378
rect 33122 37326 33124 37378
rect 33068 36932 33124 37326
rect 33180 37268 33236 38612
rect 33292 38276 33348 38286
rect 33292 38182 33348 38220
rect 33404 37490 33460 38780
rect 33852 37828 33908 39006
rect 34076 38836 34132 41020
rect 34300 41186 34468 41188
rect 34300 41134 34414 41186
rect 34466 41134 34468 41186
rect 34300 41132 34468 41134
rect 34188 40628 34244 40638
rect 34300 40628 34356 41132
rect 34412 41122 34468 41132
rect 34188 40626 34356 40628
rect 34188 40574 34190 40626
rect 34242 40574 34356 40626
rect 34188 40572 34356 40574
rect 34188 40562 34244 40572
rect 34524 40516 34580 43820
rect 34860 43876 34916 45726
rect 34972 44324 35028 44334
rect 35084 44324 35140 46396
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 35420 45892 35476 45902
rect 35532 45892 35588 46396
rect 35420 45890 35588 45892
rect 35420 45838 35422 45890
rect 35474 45838 35588 45890
rect 35420 45836 35588 45838
rect 35420 45826 35476 45836
rect 35308 45108 35364 45118
rect 35308 45014 35364 45052
rect 35532 45106 35588 45836
rect 36204 45108 36260 45118
rect 35532 45054 35534 45106
rect 35586 45054 35588 45106
rect 35532 45042 35588 45054
rect 35980 45106 36260 45108
rect 35980 45054 36206 45106
rect 36258 45054 36260 45106
rect 35980 45052 36260 45054
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 34972 44322 35084 44324
rect 34972 44270 34974 44322
rect 35026 44270 35084 44322
rect 34972 44268 35084 44270
rect 34972 44258 35028 44268
rect 35084 44230 35140 44268
rect 35868 44324 35924 44334
rect 34860 43810 34916 43820
rect 35644 44210 35700 44222
rect 35644 44158 35646 44210
rect 35698 44158 35700 44210
rect 34636 43652 34692 43662
rect 34636 43558 34692 43596
rect 34860 43538 34916 43550
rect 34860 43486 34862 43538
rect 34914 43486 34916 43538
rect 34748 43426 34804 43438
rect 34748 43374 34750 43426
rect 34802 43374 34804 43426
rect 34636 41970 34692 41982
rect 34636 41918 34638 41970
rect 34690 41918 34692 41970
rect 34636 41298 34692 41918
rect 34748 41860 34804 43374
rect 34860 43428 34916 43486
rect 34860 43362 34916 43372
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 35532 42644 35588 42654
rect 35532 42550 35588 42588
rect 35644 42308 35700 44158
rect 35756 44100 35812 44110
rect 35756 44006 35812 44044
rect 35644 42242 35700 42252
rect 34972 42196 35028 42206
rect 35028 42140 35140 42196
rect 34972 42130 35028 42140
rect 34860 42084 34916 42094
rect 34860 41990 34916 42028
rect 35084 42082 35140 42140
rect 35084 42030 35086 42082
rect 35138 42030 35140 42082
rect 35084 42018 35140 42030
rect 35644 42082 35700 42094
rect 35644 42030 35646 42082
rect 35698 42030 35700 42082
rect 35196 41972 35252 41982
rect 35196 41878 35252 41916
rect 34972 41860 35028 41870
rect 34748 41804 34916 41860
rect 34860 41412 34916 41804
rect 34972 41766 35028 41804
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 34860 41356 35028 41412
rect 34636 41246 34638 41298
rect 34690 41246 34692 41298
rect 34636 41234 34692 41246
rect 34748 41186 34804 41198
rect 34972 41188 35028 41356
rect 35644 41300 35700 42030
rect 35868 41970 35924 44268
rect 35980 44322 36036 45052
rect 36204 45042 36260 45052
rect 36428 44884 36484 44894
rect 36428 44790 36484 44828
rect 35980 44270 35982 44322
rect 36034 44270 36036 44322
rect 35980 44258 36036 44270
rect 36316 44100 36372 44110
rect 36316 44006 36372 44044
rect 36540 43652 36596 51214
rect 36652 49812 36708 49822
rect 36652 49718 36708 49756
rect 36876 49588 36932 51324
rect 36988 50932 37044 52780
rect 37100 51044 37156 56700
rect 37436 56196 37492 56206
rect 37436 56102 37492 56140
rect 37884 55412 37940 55422
rect 37884 55318 37940 55356
rect 37548 55298 37604 55310
rect 37548 55246 37550 55298
rect 37602 55246 37604 55298
rect 37212 55186 37268 55198
rect 37212 55134 37214 55186
rect 37266 55134 37268 55186
rect 37212 53956 37268 55134
rect 37324 55076 37380 55086
rect 37324 54982 37380 55020
rect 37548 55076 37604 55246
rect 38220 55300 38276 55310
rect 38220 55186 38276 55244
rect 38220 55134 38222 55186
rect 38274 55134 38276 55186
rect 37996 55076 38052 55086
rect 37548 55020 37996 55076
rect 37212 53730 37268 53900
rect 37212 53678 37214 53730
rect 37266 53678 37268 53730
rect 37212 53666 37268 53678
rect 37548 53620 37604 55020
rect 37996 54982 38052 55020
rect 38220 54740 38276 55134
rect 38220 54674 38276 54684
rect 37660 54628 37716 54638
rect 37660 54534 37716 54572
rect 38220 54516 38276 54526
rect 38220 54422 38276 54460
rect 37996 53620 38052 53630
rect 37548 53618 38052 53620
rect 37548 53566 37550 53618
rect 37602 53566 37998 53618
rect 38050 53566 38052 53618
rect 37548 53564 38052 53566
rect 37548 53554 37604 53564
rect 37212 53506 37268 53518
rect 37212 53454 37214 53506
rect 37266 53454 37268 53506
rect 37212 52162 37268 53454
rect 37212 52110 37214 52162
rect 37266 52110 37268 52162
rect 37212 52098 37268 52110
rect 37436 52274 37492 52286
rect 37436 52222 37438 52274
rect 37490 52222 37492 52274
rect 37324 51492 37380 51502
rect 37324 51378 37380 51436
rect 37324 51326 37326 51378
rect 37378 51326 37380 51378
rect 37324 51314 37380 51326
rect 37100 50978 37156 50988
rect 36988 50866 37044 50876
rect 37436 50708 37492 52222
rect 37548 51940 37604 51950
rect 37548 50818 37604 51884
rect 37548 50766 37550 50818
rect 37602 50766 37604 50818
rect 37548 50754 37604 50766
rect 37436 50642 37492 50652
rect 37324 50594 37380 50606
rect 37324 50542 37326 50594
rect 37378 50542 37380 50594
rect 37324 50428 37380 50542
rect 37660 50428 37716 53564
rect 37996 53554 38052 53564
rect 38556 53396 38612 57484
rect 40572 57428 40628 57438
rect 40460 57204 40516 57214
rect 40348 55300 40404 55310
rect 40348 55206 40404 55244
rect 38780 55076 38836 55086
rect 39116 55076 39172 55086
rect 38836 55074 39172 55076
rect 38836 55022 39118 55074
rect 39170 55022 39172 55074
rect 38836 55020 39172 55022
rect 38780 54982 38836 55020
rect 39116 55010 39172 55020
rect 39452 54514 39508 54526
rect 39452 54462 39454 54514
rect 39506 54462 39508 54514
rect 38892 54404 38948 54414
rect 38892 54310 38948 54348
rect 39004 54290 39060 54302
rect 39004 54238 39006 54290
rect 39058 54238 39060 54290
rect 39004 53732 39060 54238
rect 39004 53666 39060 53676
rect 38332 53340 38612 53396
rect 37996 53172 38052 53182
rect 37996 53078 38052 53116
rect 38332 52836 38388 53340
rect 38444 53172 38500 53182
rect 38556 53172 38612 53340
rect 39004 53508 39060 53518
rect 38892 53172 38948 53182
rect 38556 53170 38948 53172
rect 38556 53118 38894 53170
rect 38946 53118 38948 53170
rect 38556 53116 38948 53118
rect 38444 53060 38500 53116
rect 38892 53060 38948 53116
rect 38444 53004 38612 53060
rect 38444 52836 38500 52846
rect 38332 52834 38500 52836
rect 38332 52782 38446 52834
rect 38498 52782 38500 52834
rect 38332 52780 38500 52782
rect 38444 52770 38500 52780
rect 37996 52388 38052 52398
rect 36876 49522 36932 49532
rect 36988 50372 37380 50428
rect 37436 50372 37716 50428
rect 37772 51044 37828 51054
rect 36764 47012 36820 47022
rect 36988 47012 37044 50372
rect 37324 49140 37380 49150
rect 37100 49084 37324 49140
rect 37100 48466 37156 49084
rect 37324 49046 37380 49084
rect 37436 48468 37492 50372
rect 37772 49700 37828 50988
rect 37996 50818 38052 52332
rect 38556 52276 38612 53004
rect 38892 52994 38948 53004
rect 39004 52948 39060 53452
rect 39452 53284 39508 54462
rect 39788 54516 39844 54526
rect 39788 54422 39844 54460
rect 39564 54404 39620 54414
rect 39564 54310 39620 54348
rect 39788 53956 39844 53966
rect 39676 53730 39732 53742
rect 39676 53678 39678 53730
rect 39730 53678 39732 53730
rect 39676 53508 39732 53678
rect 39676 53442 39732 53452
rect 39340 53228 39508 53284
rect 39004 52882 39060 52892
rect 39228 53060 39284 53070
rect 39004 52276 39060 52286
rect 38556 52274 39060 52276
rect 38556 52222 38558 52274
rect 38610 52222 39006 52274
rect 39058 52222 39060 52274
rect 38556 52220 39060 52222
rect 38556 52182 38612 52220
rect 39004 52210 39060 52220
rect 38108 52050 38164 52062
rect 38108 51998 38110 52050
rect 38162 51998 38164 52050
rect 38108 51492 38164 51998
rect 38444 51940 38500 51950
rect 38444 51846 38500 51884
rect 38108 51426 38164 51436
rect 38444 51490 38500 51502
rect 38444 51438 38446 51490
rect 38498 51438 38500 51490
rect 37996 50766 37998 50818
rect 38050 50766 38052 50818
rect 37996 50754 38052 50766
rect 38108 50820 38164 50830
rect 38108 50726 38164 50764
rect 38332 50708 38388 50718
rect 38444 50708 38500 51438
rect 38388 50652 38500 50708
rect 39228 50706 39284 53004
rect 39228 50654 39230 50706
rect 39282 50654 39284 50706
rect 38332 50642 38388 50652
rect 39228 50642 39284 50654
rect 37996 50596 38052 50606
rect 37996 50502 38052 50540
rect 38780 50484 38836 50494
rect 39340 50428 39396 53228
rect 39564 53172 39620 53182
rect 39564 53078 39620 53116
rect 39788 53170 39844 53900
rect 40012 53844 40068 53854
rect 40012 53750 40068 53788
rect 40348 53620 40404 53630
rect 40348 53526 40404 53564
rect 39788 53118 39790 53170
rect 39842 53118 39844 53170
rect 39788 53106 39844 53118
rect 40124 53172 40180 53182
rect 39452 53060 39508 53070
rect 39452 52966 39508 53004
rect 40012 53060 40068 53070
rect 39452 52276 39508 52286
rect 39452 52164 39508 52220
rect 39452 52162 39620 52164
rect 39452 52110 39454 52162
rect 39506 52110 39620 52162
rect 39452 52108 39620 52110
rect 39452 52098 39508 52108
rect 39564 51492 39620 52108
rect 40012 52162 40068 53004
rect 40012 52110 40014 52162
rect 40066 52110 40068 52162
rect 39676 51940 39732 51950
rect 39676 51846 39732 51884
rect 39900 51604 39956 51614
rect 40012 51604 40068 52110
rect 39900 51602 40068 51604
rect 39900 51550 39902 51602
rect 39954 51550 40068 51602
rect 39900 51548 40068 51550
rect 40124 52050 40180 53116
rect 40124 51998 40126 52050
rect 40178 51998 40180 52050
rect 40124 51602 40180 51998
rect 40124 51550 40126 51602
rect 40178 51550 40180 51602
rect 39900 51538 39956 51548
rect 39676 51492 39732 51502
rect 39564 51490 39732 51492
rect 39564 51438 39678 51490
rect 39730 51438 39732 51490
rect 39564 51436 39732 51438
rect 39676 51426 39732 51436
rect 40124 51268 40180 51550
rect 39676 51212 40180 51268
rect 40236 52164 40292 52174
rect 39564 50708 39620 50718
rect 38780 50372 38948 50428
rect 39340 50372 39508 50428
rect 38444 50036 38500 50046
rect 37996 49700 38052 49710
rect 37772 49698 38164 49700
rect 37772 49646 37998 49698
rect 38050 49646 38164 49698
rect 37772 49644 38164 49646
rect 37996 49634 38052 49644
rect 37996 49140 38052 49150
rect 37100 48414 37102 48466
rect 37154 48414 37156 48466
rect 37100 48132 37156 48414
rect 37100 48066 37156 48076
rect 37324 48412 37492 48468
rect 37548 49026 37604 49038
rect 37548 48974 37550 49026
rect 37602 48974 37604 49026
rect 37212 47460 37268 47470
rect 37212 47366 37268 47404
rect 36988 46956 37156 47012
rect 36652 46562 36708 46574
rect 36652 46510 36654 46562
rect 36706 46510 36708 46562
rect 36652 45780 36708 46510
rect 36764 46562 36820 46956
rect 36764 46510 36766 46562
rect 36818 46510 36820 46562
rect 36764 46498 36820 46510
rect 36988 46674 37044 46686
rect 36988 46622 36990 46674
rect 37042 46622 37044 46674
rect 36988 46564 37044 46622
rect 36652 45714 36708 45724
rect 36876 45556 36932 45566
rect 36764 44212 36820 44222
rect 36652 43652 36708 43662
rect 36540 43650 36708 43652
rect 36540 43598 36654 43650
rect 36706 43598 36708 43650
rect 36540 43596 36708 43598
rect 36428 43540 36484 43550
rect 36428 43446 36484 43484
rect 36316 42980 36372 42990
rect 36316 42886 36372 42924
rect 35868 41918 35870 41970
rect 35922 41918 35924 41970
rect 35868 41906 35924 41918
rect 36092 42754 36148 42766
rect 36092 42702 36094 42754
rect 36146 42702 36148 42754
rect 34748 41134 34750 41186
rect 34802 41134 34804 41186
rect 34748 41076 34804 41134
rect 34748 41010 34804 41020
rect 34860 41132 35028 41188
rect 35084 41244 35700 41300
rect 35084 41186 35140 41244
rect 35084 41134 35086 41186
rect 35138 41134 35140 41186
rect 34860 40626 34916 41132
rect 35084 40628 35140 41134
rect 34860 40574 34862 40626
rect 34914 40574 34916 40626
rect 34860 40562 34916 40574
rect 34972 40572 35140 40628
rect 34300 40460 34580 40516
rect 34972 40514 35028 40572
rect 34972 40462 34974 40514
rect 35026 40462 35028 40514
rect 34300 39618 34356 40460
rect 34972 40450 35028 40462
rect 35084 40404 35140 40414
rect 35084 40310 35140 40348
rect 35196 40402 35252 40414
rect 35196 40350 35198 40402
rect 35250 40350 35252 40402
rect 35196 40180 35252 40350
rect 34748 40124 35252 40180
rect 35308 40180 35364 41244
rect 35420 40404 35476 40414
rect 35420 40402 35924 40404
rect 35420 40350 35422 40402
rect 35474 40350 35924 40402
rect 35420 40348 35924 40350
rect 35420 40338 35476 40348
rect 35308 40124 35588 40180
rect 34300 39566 34302 39618
rect 34354 39566 34356 39618
rect 34300 39396 34356 39566
rect 34300 39330 34356 39340
rect 34412 39620 34468 39630
rect 34188 38836 34244 38846
rect 34076 38780 34188 38836
rect 34244 38780 34356 38836
rect 34188 38770 34244 38780
rect 34300 38500 34356 38780
rect 34412 38724 34468 39564
rect 34412 38612 34580 38668
rect 34300 38444 34468 38500
rect 34188 38164 34244 38174
rect 34188 38070 34244 38108
rect 34300 37828 34356 37838
rect 33852 37772 34132 37828
rect 33404 37438 33406 37490
rect 33458 37438 33460 37490
rect 33404 37426 33460 37438
rect 33516 37604 33572 37614
rect 33180 37202 33236 37212
rect 33124 36876 33348 36932
rect 33068 36866 33124 36876
rect 33012 36652 33236 36708
rect 32956 36614 33012 36652
rect 32620 36318 32622 36370
rect 32674 36318 32676 36370
rect 32620 36306 32676 36318
rect 33180 36370 33236 36652
rect 33292 36482 33348 36876
rect 33516 36594 33572 37548
rect 34076 37378 34132 37772
rect 34300 37734 34356 37772
rect 34076 37326 34078 37378
rect 34130 37326 34132 37378
rect 34076 37314 34132 37326
rect 33964 37268 34020 37278
rect 33516 36542 33518 36594
rect 33570 36542 33572 36594
rect 33516 36530 33572 36542
rect 33852 37266 34020 37268
rect 33852 37214 33966 37266
rect 34018 37214 34020 37266
rect 33852 37212 34020 37214
rect 33292 36430 33294 36482
rect 33346 36430 33348 36482
rect 33292 36418 33348 36430
rect 33180 36318 33182 36370
rect 33234 36318 33236 36370
rect 33180 36306 33236 36318
rect 33852 36148 33908 37212
rect 33964 37202 34020 37212
rect 33964 36484 34020 36494
rect 33964 36390 34020 36428
rect 34076 36372 34132 36382
rect 34076 36278 34132 36316
rect 34412 36370 34468 38444
rect 34524 38050 34580 38612
rect 34524 37998 34526 38050
rect 34578 37998 34580 38050
rect 34524 37986 34580 37998
rect 34748 36820 34804 40124
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 34860 39620 34916 39630
rect 35420 39620 35476 39630
rect 35532 39620 35588 40124
rect 35868 39730 35924 40348
rect 35868 39678 35870 39730
rect 35922 39678 35924 39730
rect 35868 39666 35924 39678
rect 36092 39732 36148 42702
rect 36652 42644 36708 43596
rect 36764 43650 36820 44156
rect 36764 43598 36766 43650
rect 36818 43598 36820 43650
rect 36764 43586 36820 43598
rect 36652 42578 36708 42588
rect 36652 42308 36708 42318
rect 36540 40964 36596 40974
rect 36148 39676 36484 39732
rect 36092 39666 36148 39676
rect 34860 39526 34916 39564
rect 35196 39618 35588 39620
rect 35196 39566 35422 39618
rect 35474 39566 35588 39618
rect 35196 39564 35588 39566
rect 35196 39058 35252 39564
rect 35420 39554 35476 39564
rect 35756 39508 35812 39518
rect 35756 39414 35812 39452
rect 35980 39396 36036 39406
rect 35980 39302 36036 39340
rect 35196 39006 35198 39058
rect 35250 39006 35252 39058
rect 35196 38994 35252 39006
rect 36316 39060 36372 39070
rect 34860 38948 34916 38958
rect 34860 38668 34916 38892
rect 35756 38948 35812 38958
rect 35756 38854 35812 38892
rect 35532 38834 35588 38846
rect 35532 38782 35534 38834
rect 35586 38782 35588 38834
rect 34860 38612 35028 38668
rect 34860 38050 34916 38062
rect 34860 37998 34862 38050
rect 34914 37998 34916 38050
rect 34860 37380 34916 37998
rect 34860 37314 34916 37324
rect 34972 37938 35028 38612
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 34972 37886 34974 37938
rect 35026 37886 35028 37938
rect 34412 36318 34414 36370
rect 34466 36318 34468 36370
rect 34412 36306 34468 36318
rect 34524 36764 34804 36820
rect 32508 36092 33124 36148
rect 32508 35586 32564 35598
rect 32508 35534 32510 35586
rect 32562 35534 32564 35586
rect 32508 35476 32564 35534
rect 32508 35410 32564 35420
rect 33068 35140 33124 36092
rect 33852 36082 33908 36092
rect 34188 36258 34244 36270
rect 34188 36206 34190 36258
rect 34242 36206 34244 36258
rect 33180 35698 33236 35710
rect 33180 35646 33182 35698
rect 33234 35646 33236 35698
rect 33180 35476 33236 35646
rect 33180 35410 33236 35420
rect 33628 35698 33684 35710
rect 33628 35646 33630 35698
rect 33682 35646 33684 35698
rect 33292 35140 33348 35150
rect 32284 35084 32452 35140
rect 33068 35138 33348 35140
rect 33068 35086 33294 35138
rect 33346 35086 33348 35138
rect 33068 35084 33348 35086
rect 32284 34916 32340 34926
rect 32172 34914 32340 34916
rect 32172 34862 32286 34914
rect 32338 34862 32340 34914
rect 32172 34860 32340 34862
rect 32284 34850 32340 34860
rect 32060 34638 32062 34690
rect 32114 34638 32116 34690
rect 32060 34356 32116 34638
rect 32060 34290 32116 34300
rect 31052 33966 31054 34018
rect 31106 33966 31108 34018
rect 28588 33122 28644 33134
rect 28588 33070 28590 33122
rect 28642 33070 28644 33122
rect 28588 32788 28644 33070
rect 29484 33122 29540 33134
rect 29484 33070 29486 33122
rect 29538 33070 29540 33122
rect 28588 32722 28644 32732
rect 29260 32786 29316 32798
rect 29260 32734 29262 32786
rect 29314 32734 29316 32786
rect 29260 32452 29316 32734
rect 29484 32788 29540 33070
rect 29820 33124 29876 33134
rect 30268 33124 30324 33134
rect 29820 33122 30324 33124
rect 29820 33070 29822 33122
rect 29874 33070 30270 33122
rect 30322 33070 30324 33122
rect 29820 33068 30324 33070
rect 29820 33058 29876 33068
rect 29484 32722 29540 32732
rect 29820 32788 29876 32798
rect 29820 32694 29876 32732
rect 30156 32564 30212 32574
rect 30268 32564 30324 33068
rect 30212 32508 30324 32564
rect 30156 32470 30212 32508
rect 29260 32386 29316 32396
rect 28476 31714 28532 31724
rect 30044 31778 30100 31790
rect 30044 31726 30046 31778
rect 30098 31726 30100 31778
rect 25900 31502 25902 31554
rect 25954 31502 25956 31554
rect 25564 30994 25620 31006
rect 25564 30942 25566 30994
rect 25618 30942 25620 30994
rect 25564 30884 25620 30942
rect 25564 30818 25620 30828
rect 25900 30884 25956 31502
rect 28140 31332 28196 31342
rect 26908 30996 26964 31006
rect 26908 30902 26964 30940
rect 25900 30818 25956 30828
rect 26236 30884 26292 30894
rect 26236 30790 26292 30828
rect 27804 30324 27860 30334
rect 25004 30158 25006 30210
rect 25058 30158 25060 30210
rect 25004 30146 25060 30158
rect 25340 30210 25396 30222
rect 25340 30158 25342 30210
rect 25394 30158 25396 30210
rect 24668 29598 24670 29650
rect 24722 29598 24724 29650
rect 24668 29540 24724 29598
rect 25116 29652 25172 29662
rect 25172 29596 25284 29652
rect 25116 29586 25172 29596
rect 24668 29474 24724 29484
rect 25228 29538 25284 29596
rect 25340 29650 25396 30158
rect 25340 29598 25342 29650
rect 25394 29598 25396 29650
rect 25340 29586 25396 29598
rect 25676 29988 25732 29998
rect 25228 29486 25230 29538
rect 25282 29486 25284 29538
rect 25228 29474 25284 29486
rect 25452 29540 25508 29550
rect 25452 29426 25508 29484
rect 25452 29374 25454 29426
rect 25506 29374 25508 29426
rect 25452 29362 25508 29374
rect 25676 29426 25732 29932
rect 26236 29540 26292 29550
rect 26236 29446 26292 29484
rect 25676 29374 25678 29426
rect 25730 29374 25732 29426
rect 25676 29362 25732 29374
rect 24444 29150 24446 29202
rect 24498 29150 24500 29202
rect 24444 29138 24500 29150
rect 24780 29202 24836 29214
rect 24780 29150 24782 29202
rect 24834 29150 24836 29202
rect 24220 28756 24276 28766
rect 24108 28754 24612 28756
rect 24108 28702 24222 28754
rect 24274 28702 24612 28754
rect 24108 28700 24612 28702
rect 24220 28690 24276 28700
rect 22540 27794 22596 27804
rect 22652 28588 22764 28644
rect 22820 28588 22932 28644
rect 24556 28642 24612 28700
rect 24556 28590 24558 28642
rect 24610 28590 24612 28642
rect 22316 27186 22484 27188
rect 22316 27134 22318 27186
rect 22370 27134 22484 27186
rect 22316 27132 22484 27134
rect 22316 27122 22372 27132
rect 21756 26852 22260 26908
rect 21588 25340 21700 25396
rect 21756 26292 21812 26302
rect 21756 25618 21812 26236
rect 22204 26290 22260 26852
rect 22204 26238 22206 26290
rect 22258 26238 22260 26290
rect 22204 25956 22260 26238
rect 22204 25890 22260 25900
rect 21756 25566 21758 25618
rect 21810 25566 21812 25618
rect 20748 24052 20804 24062
rect 20636 23996 20748 24052
rect 20748 23958 20804 23996
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19628 23102 19630 23154
rect 19682 23102 19684 23154
rect 19628 23090 19684 23102
rect 20300 23156 20356 23166
rect 20188 22820 20244 22830
rect 19740 22372 19796 22382
rect 19740 22278 19796 22316
rect 20188 22372 20244 22764
rect 20300 22482 20356 23100
rect 20300 22430 20302 22482
rect 20354 22430 20356 22482
rect 20300 22418 20356 22430
rect 20636 23154 20692 23166
rect 20636 23102 20638 23154
rect 20690 23102 20692 23154
rect 20188 22306 20244 22316
rect 20412 22372 20468 22382
rect 20188 22148 20244 22158
rect 19404 22092 19572 22148
rect 19292 20690 19348 21420
rect 19404 20804 19460 20814
rect 19404 20710 19460 20748
rect 19292 20638 19294 20690
rect 19346 20638 19348 20690
rect 19292 20580 19348 20638
rect 19292 20524 19460 20580
rect 19404 20468 19460 20524
rect 19180 20412 19348 20468
rect 19068 19170 19124 19180
rect 19180 20244 19236 20254
rect 19180 20130 19236 20188
rect 19180 20078 19182 20130
rect 19234 20078 19236 20130
rect 19180 19234 19236 20078
rect 19292 19796 19348 20412
rect 19404 20402 19460 20412
rect 19292 19730 19348 19740
rect 19404 20018 19460 20030
rect 19404 19966 19406 20018
rect 19458 19966 19460 20018
rect 19180 19182 19182 19234
rect 19234 19182 19236 19234
rect 19180 19170 19236 19182
rect 19292 19236 19348 19246
rect 19404 19236 19460 19966
rect 19348 19180 19460 19236
rect 19292 19170 19348 19180
rect 19180 19012 19236 19022
rect 19068 18116 19124 18126
rect 19068 17666 19124 18060
rect 19068 17614 19070 17666
rect 19122 17614 19124 17666
rect 19068 17602 19124 17614
rect 19180 17444 19236 18956
rect 19404 18676 19460 18686
rect 19404 18582 19460 18620
rect 19292 17780 19348 17790
rect 19292 17666 19348 17724
rect 19292 17614 19294 17666
rect 19346 17614 19348 17666
rect 19292 17602 19348 17614
rect 19180 17388 19348 17444
rect 18956 17276 19124 17332
rect 18844 16882 18900 16894
rect 18844 16830 18846 16882
rect 18898 16830 18900 16882
rect 18844 16324 18900 16830
rect 18844 16258 18900 16268
rect 18732 15222 18788 15260
rect 18956 15202 19012 15214
rect 18956 15150 18958 15202
rect 19010 15150 19012 15202
rect 18732 14420 18788 14430
rect 18508 14418 18788 14420
rect 18508 14366 18734 14418
rect 18786 14366 18788 14418
rect 18508 14364 18788 14366
rect 18732 14354 18788 14364
rect 18396 14140 18900 14196
rect 18396 13636 18452 13646
rect 17836 13186 18004 13188
rect 17836 13134 17838 13186
rect 17890 13134 18004 13186
rect 17836 13132 18004 13134
rect 18284 13580 18396 13636
rect 17836 13122 17892 13132
rect 17612 13076 17668 13086
rect 17388 12798 17390 12850
rect 17442 12798 17444 12850
rect 17388 11620 17444 12798
rect 17500 13074 17668 13076
rect 17500 13022 17614 13074
rect 17666 13022 17668 13074
rect 17500 13020 17668 13022
rect 17500 12404 17556 13020
rect 17612 13010 17668 13020
rect 17500 12338 17556 12348
rect 17612 12852 17668 12862
rect 17500 12066 17556 12078
rect 17500 12014 17502 12066
rect 17554 12014 17556 12066
rect 17500 11844 17556 12014
rect 17500 11778 17556 11788
rect 17388 11564 17556 11620
rect 17388 11396 17444 11406
rect 17388 11302 17444 11340
rect 17276 9996 17444 10052
rect 17276 9826 17332 9838
rect 17276 9774 17278 9826
rect 17330 9774 17332 9826
rect 17276 9604 17332 9774
rect 17276 9538 17332 9548
rect 17052 9100 17220 9156
rect 16828 9044 16884 9054
rect 16828 8484 16884 8988
rect 16940 9044 16996 9054
rect 17052 9044 17108 9100
rect 16940 9042 17108 9044
rect 16940 8990 16942 9042
rect 16994 8990 17108 9042
rect 16940 8988 17108 8990
rect 16940 8978 16996 8988
rect 17164 8708 17220 9100
rect 17164 8642 17220 8652
rect 16828 8428 17108 8484
rect 16716 8306 16772 8316
rect 16828 8260 16884 8270
rect 16828 8166 16884 8204
rect 16604 7980 16996 8036
rect 16940 7698 16996 7980
rect 16940 7646 16942 7698
rect 16994 7646 16996 7698
rect 16940 7634 16996 7646
rect 16492 6860 16772 6916
rect 16156 6750 16158 6802
rect 16210 6750 16212 6802
rect 16156 6738 16212 6750
rect 16044 6244 16100 6636
rect 16604 6690 16660 6702
rect 16604 6638 16606 6690
rect 16658 6638 16660 6690
rect 16492 6580 16548 6590
rect 16380 6524 16492 6580
rect 16044 6188 16324 6244
rect 16268 5908 16324 6188
rect 16268 5814 16324 5852
rect 16156 5796 16212 5806
rect 15708 5794 16212 5796
rect 15708 5742 16158 5794
rect 16210 5742 16212 5794
rect 15708 5740 16212 5742
rect 16156 5730 16212 5740
rect 15484 5122 15652 5124
rect 15484 5070 15486 5122
rect 15538 5070 15652 5122
rect 15484 5068 15652 5070
rect 15708 5572 15764 5582
rect 15484 5058 15540 5068
rect 15036 4956 15316 5012
rect 14924 4900 14980 4910
rect 14924 4806 14980 4844
rect 15260 4676 15316 4686
rect 15260 4562 15316 4620
rect 15596 4564 15652 4574
rect 15708 4564 15764 5516
rect 16268 5236 16324 5246
rect 16380 5236 16436 6524
rect 16492 6514 16548 6524
rect 16604 5796 16660 6638
rect 16268 5234 16436 5236
rect 16268 5182 16270 5234
rect 16322 5182 16436 5234
rect 16268 5180 16436 5182
rect 16268 5170 16324 5180
rect 15260 4510 15262 4562
rect 15314 4510 15316 4562
rect 15260 4498 15316 4510
rect 15372 4562 15764 4564
rect 15372 4510 15598 4562
rect 15650 4510 15764 4562
rect 15372 4508 15764 4510
rect 15820 5010 15876 5022
rect 15820 4958 15822 5010
rect 15874 4958 15876 5010
rect 15820 4900 15876 4958
rect 14924 3668 14980 3678
rect 14812 3666 14980 3668
rect 14812 3614 14926 3666
rect 14978 3614 14980 3666
rect 14812 3612 14980 3614
rect 14924 3602 14980 3612
rect 15372 3666 15428 4508
rect 15596 4498 15652 4508
rect 15820 4228 15876 4844
rect 16380 4900 16436 5180
rect 16380 4834 16436 4844
rect 16492 5682 16548 5694
rect 16492 5630 16494 5682
rect 16546 5630 16548 5682
rect 16492 4564 16548 5630
rect 16604 5460 16660 5740
rect 16604 5394 16660 5404
rect 16716 5460 16772 6860
rect 16940 6132 16996 6142
rect 16828 5460 16884 5470
rect 16716 5404 16828 5460
rect 16604 5124 16660 5134
rect 16604 5010 16660 5068
rect 16604 4958 16606 5010
rect 16658 4958 16660 5010
rect 16604 4946 16660 4958
rect 16492 4508 16660 4564
rect 15820 4162 15876 4172
rect 16492 4226 16548 4238
rect 16492 4174 16494 4226
rect 16546 4174 16548 4226
rect 16492 4114 16548 4174
rect 16492 4062 16494 4114
rect 16546 4062 16548 4114
rect 16492 4050 16548 4062
rect 16492 3892 16548 3902
rect 15372 3614 15374 3666
rect 15426 3614 15428 3666
rect 15372 3602 15428 3614
rect 15820 3668 15876 3678
rect 15820 3574 15876 3612
rect 16492 3666 16548 3836
rect 16492 3614 16494 3666
rect 16546 3614 16548 3666
rect 16492 3602 16548 3614
rect 13244 2706 13300 2716
rect 16604 2660 16660 4508
rect 16716 4114 16772 5404
rect 16828 5394 16884 5404
rect 16940 5122 16996 6076
rect 16940 5070 16942 5122
rect 16994 5070 16996 5122
rect 16940 5058 16996 5070
rect 16716 4062 16718 4114
rect 16770 4062 16772 4114
rect 16716 4050 16772 4062
rect 16940 4900 16996 4910
rect 16940 4562 16996 4844
rect 16940 4510 16942 4562
rect 16994 4510 16996 4562
rect 16940 4004 16996 4510
rect 16940 3938 16996 3948
rect 17052 3778 17108 8428
rect 17388 8372 17444 9996
rect 17500 9156 17556 11564
rect 17612 10834 17668 12796
rect 17612 10782 17614 10834
rect 17666 10782 17668 10834
rect 17612 10770 17668 10782
rect 17836 12404 17892 12414
rect 17836 10500 17892 12348
rect 17948 12290 18004 12302
rect 17948 12238 17950 12290
rect 18002 12238 18004 12290
rect 17948 10834 18004 12238
rect 18172 12178 18228 12190
rect 18172 12126 18174 12178
rect 18226 12126 18228 12178
rect 18172 11284 18228 12126
rect 18172 11218 18228 11228
rect 17948 10782 17950 10834
rect 18002 10782 18004 10834
rect 17948 10770 18004 10782
rect 18172 10836 18228 10846
rect 18060 10724 18116 10734
rect 18060 10610 18116 10668
rect 18060 10558 18062 10610
rect 18114 10558 18116 10610
rect 18060 10546 18116 10558
rect 17948 10500 18004 10510
rect 17836 10498 18004 10500
rect 17836 10446 17950 10498
rect 18002 10446 18004 10498
rect 17836 10444 18004 10446
rect 17948 9268 18004 10444
rect 18060 10388 18116 10398
rect 18060 9828 18116 10332
rect 18060 9380 18116 9772
rect 18172 9826 18228 10780
rect 18172 9774 18174 9826
rect 18226 9774 18228 9826
rect 18172 9604 18228 9774
rect 18172 9538 18228 9548
rect 18060 9324 18228 9380
rect 17948 9212 18116 9268
rect 17500 9100 17892 9156
rect 17276 8316 17444 8372
rect 17500 8818 17556 8830
rect 17500 8766 17502 8818
rect 17554 8766 17556 8818
rect 17276 5908 17332 8316
rect 17276 5684 17332 5852
rect 17276 5618 17332 5628
rect 17388 8148 17444 8158
rect 17388 5572 17444 8092
rect 17500 8146 17556 8766
rect 17612 8708 17668 8718
rect 17668 8652 17780 8708
rect 17612 8642 17668 8652
rect 17500 8094 17502 8146
rect 17554 8094 17556 8146
rect 17500 8082 17556 8094
rect 17388 5124 17444 5516
rect 17612 7588 17668 7598
rect 17612 5460 17668 7532
rect 17724 6018 17780 8652
rect 17836 7698 17892 9100
rect 17836 7646 17838 7698
rect 17890 7646 17892 7698
rect 17836 6132 17892 7646
rect 17948 9042 18004 9054
rect 17948 8990 17950 9042
rect 18002 8990 18004 9042
rect 17948 7700 18004 8990
rect 17948 7634 18004 7644
rect 17948 7476 18004 7486
rect 17948 7362 18004 7420
rect 17948 7310 17950 7362
rect 18002 7310 18004 7362
rect 17948 7298 18004 7310
rect 18060 6804 18116 9212
rect 18172 9042 18228 9324
rect 18172 8990 18174 9042
rect 18226 8990 18228 9042
rect 18172 8820 18228 8990
rect 18172 8754 18228 8764
rect 18284 8484 18340 13580
rect 18396 13542 18452 13580
rect 18508 13524 18564 13534
rect 18396 11508 18452 11518
rect 18396 11414 18452 11452
rect 18508 11508 18564 13468
rect 18844 12962 18900 14140
rect 18956 13748 19012 15150
rect 18956 13524 19012 13692
rect 18956 13458 19012 13468
rect 18844 12910 18846 12962
rect 18898 12910 18900 12962
rect 18844 11788 18900 12910
rect 18956 13186 19012 13198
rect 18956 13134 18958 13186
rect 19010 13134 19012 13186
rect 18956 12180 19012 13134
rect 18956 12114 19012 12124
rect 18732 11732 18900 11788
rect 18956 11956 19012 11966
rect 18620 11508 18676 11518
rect 18508 11452 18620 11508
rect 18508 10948 18564 11452
rect 18620 11442 18676 11452
rect 18508 10882 18564 10892
rect 18396 10500 18452 10510
rect 18396 9716 18452 10444
rect 18620 9828 18676 9838
rect 18396 9650 18452 9660
rect 18508 9772 18620 9828
rect 18396 9492 18452 9502
rect 18396 8708 18452 9436
rect 18508 9154 18564 9772
rect 18620 9762 18676 9772
rect 18508 9102 18510 9154
rect 18562 9102 18564 9154
rect 18508 9090 18564 9102
rect 18620 9604 18676 9614
rect 18396 8642 18452 8652
rect 18508 8596 18564 8606
rect 18284 8428 18452 8484
rect 18172 8260 18228 8270
rect 18172 7924 18228 8204
rect 18172 6914 18228 7868
rect 18172 6862 18174 6914
rect 18226 6862 18228 6914
rect 18172 6850 18228 6862
rect 18396 8148 18452 8428
rect 18508 8258 18564 8540
rect 18508 8206 18510 8258
rect 18562 8206 18564 8258
rect 18508 8194 18564 8206
rect 18060 6692 18116 6748
rect 18284 6804 18340 6814
rect 18060 6636 18228 6692
rect 17836 6066 17892 6076
rect 17724 5966 17726 6018
rect 17778 5966 17780 6018
rect 17724 5954 17780 5966
rect 17836 5906 17892 5918
rect 17836 5854 17838 5906
rect 17890 5854 17892 5906
rect 17612 5404 17780 5460
rect 17612 5124 17668 5134
rect 17388 5122 17668 5124
rect 17388 5070 17614 5122
rect 17666 5070 17668 5122
rect 17388 5068 17668 5070
rect 17612 5058 17668 5068
rect 17052 3726 17054 3778
rect 17106 3726 17108 3778
rect 17052 3714 17108 3726
rect 17276 4900 17332 4910
rect 17276 3666 17332 4844
rect 17612 4564 17668 4574
rect 17612 4470 17668 4508
rect 17276 3614 17278 3666
rect 17330 3614 17332 3666
rect 17276 3602 17332 3614
rect 17724 3666 17780 5404
rect 17836 5124 17892 5854
rect 18060 5796 18116 5806
rect 17836 5030 17892 5068
rect 17948 5124 18004 5134
rect 18060 5124 18116 5740
rect 17948 5122 18116 5124
rect 17948 5070 17950 5122
rect 18002 5070 18116 5122
rect 17948 5068 18116 5070
rect 17948 5058 18004 5068
rect 18172 4452 18228 6636
rect 18284 5906 18340 6748
rect 18396 6692 18452 8092
rect 18620 7700 18676 9548
rect 18732 9380 18788 11732
rect 18956 11394 19012 11900
rect 18956 11342 18958 11394
rect 19010 11342 19012 11394
rect 18956 11330 19012 11342
rect 19068 10836 19124 17276
rect 19180 16548 19236 16558
rect 19180 15426 19236 16492
rect 19180 15374 19182 15426
rect 19234 15374 19236 15426
rect 19180 15362 19236 15374
rect 19292 15428 19348 17388
rect 19516 16882 19572 22092
rect 19628 22036 19684 22046
rect 19628 20132 19684 21980
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19964 21812 20020 21822
rect 19852 21474 19908 21486
rect 19852 21422 19854 21474
rect 19906 21422 19908 21474
rect 19852 20580 19908 21422
rect 19964 21252 20020 21756
rect 20188 21698 20244 22092
rect 20188 21646 20190 21698
rect 20242 21646 20244 21698
rect 20188 21634 20244 21646
rect 20300 21588 20356 21598
rect 20300 21494 20356 21532
rect 20412 21364 20468 22316
rect 19964 21186 20020 21196
rect 20300 21308 20468 21364
rect 19852 20514 19908 20524
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19740 20132 19796 20142
rect 19628 20130 19796 20132
rect 19628 20078 19742 20130
rect 19794 20078 19796 20130
rect 19628 20076 19796 20078
rect 19740 20066 19796 20076
rect 20076 20018 20132 20030
rect 20076 19966 20078 20018
rect 20130 19966 20132 20018
rect 20076 19796 20132 19966
rect 20076 19730 20132 19740
rect 20300 19234 20356 21308
rect 20636 20804 20692 23102
rect 20748 22484 20804 22494
rect 20748 22390 20804 22428
rect 20860 22260 20916 25340
rect 21532 25302 21588 25340
rect 21756 25284 21812 25566
rect 22316 25508 22372 25518
rect 22316 25414 22372 25452
rect 21756 25218 21812 25228
rect 22316 24948 22372 24958
rect 20972 24836 21028 24846
rect 20972 24742 21028 24780
rect 21420 24836 21476 24846
rect 21196 24610 21252 24622
rect 21196 24558 21198 24610
rect 21250 24558 21252 24610
rect 20636 20738 20692 20748
rect 20748 22204 20916 22260
rect 20972 22596 21028 22606
rect 20412 20580 20468 20590
rect 20412 20132 20468 20524
rect 20636 20580 20692 20590
rect 20636 20486 20692 20524
rect 20468 20076 20580 20132
rect 20412 20066 20468 20076
rect 20300 19182 20302 19234
rect 20354 19182 20356 19234
rect 20300 19170 20356 19182
rect 20412 19906 20468 19918
rect 20412 19854 20414 19906
rect 20466 19854 20468 19906
rect 20412 19236 20468 19854
rect 20412 19170 20468 19180
rect 19964 19122 20020 19134
rect 19964 19070 19966 19122
rect 20018 19070 20020 19122
rect 19964 19012 20020 19070
rect 19628 18956 20020 19012
rect 20412 19012 20468 19022
rect 19628 18452 19684 18956
rect 20412 18918 20468 18956
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19628 17780 19684 18396
rect 20076 18452 20132 18462
rect 20076 18450 20244 18452
rect 20076 18398 20078 18450
rect 20130 18398 20244 18450
rect 20076 18396 20244 18398
rect 20076 18386 20132 18396
rect 20188 18116 20244 18396
rect 20188 18050 20244 18060
rect 19628 17714 19684 17724
rect 20412 17892 20468 17902
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19516 16830 19518 16882
rect 19570 16830 19572 16882
rect 19516 16818 19572 16830
rect 19292 15362 19348 15372
rect 19404 16772 19460 16782
rect 19292 14308 19348 14318
rect 19180 13860 19236 13870
rect 19180 13746 19236 13804
rect 19180 13694 19182 13746
rect 19234 13694 19236 13746
rect 19180 11844 19236 13694
rect 19180 11778 19236 11788
rect 19068 10770 19124 10780
rect 18956 10612 19012 10622
rect 18956 10518 19012 10556
rect 19292 10164 19348 14252
rect 19404 13634 19460 16716
rect 19852 16660 19908 16670
rect 19852 16566 19908 16604
rect 19964 16324 20020 16334
rect 19852 16268 19964 16324
rect 19740 16212 19796 16222
rect 19740 16118 19796 16156
rect 19852 15988 19908 16268
rect 19964 16258 20020 16268
rect 19964 16100 20020 16110
rect 20188 16100 20244 16110
rect 19964 16098 20244 16100
rect 19964 16046 19966 16098
rect 20018 16046 20190 16098
rect 20242 16046 20244 16098
rect 19964 16044 20244 16046
rect 19964 16034 20020 16044
rect 20188 16034 20244 16044
rect 19516 15986 19908 15988
rect 19516 15934 19854 15986
rect 19906 15934 19908 15986
rect 19516 15932 19908 15934
rect 19516 14084 19572 15932
rect 19852 15922 19908 15932
rect 20412 15986 20468 17836
rect 20524 16772 20580 20076
rect 20636 17442 20692 17454
rect 20636 17390 20638 17442
rect 20690 17390 20692 17442
rect 20636 17332 20692 17390
rect 20636 16994 20692 17276
rect 20636 16942 20638 16994
rect 20690 16942 20692 16994
rect 20636 16930 20692 16942
rect 20524 16716 20692 16772
rect 20412 15934 20414 15986
rect 20466 15934 20468 15986
rect 20412 15922 20468 15934
rect 20524 16436 20580 16446
rect 20524 16098 20580 16380
rect 20524 16046 20526 16098
rect 20578 16046 20580 16098
rect 20524 15876 20580 16046
rect 20524 15810 20580 15820
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20636 15652 20692 16716
rect 19836 15642 20100 15652
rect 20524 15596 20692 15652
rect 19516 14018 19572 14028
rect 19628 15540 19684 15550
rect 19404 13582 19406 13634
rect 19458 13582 19460 13634
rect 19404 13570 19460 13582
rect 19404 12962 19460 12974
rect 19404 12910 19406 12962
rect 19458 12910 19460 12962
rect 19404 10724 19460 12910
rect 19628 12404 19684 15484
rect 19740 15428 19796 15438
rect 19740 14308 19796 15372
rect 20300 15314 20356 15326
rect 20300 15262 20302 15314
rect 20354 15262 20356 15314
rect 20188 15202 20244 15214
rect 20188 15150 20190 15202
rect 20242 15150 20244 15202
rect 20188 15092 20244 15150
rect 20188 15026 20244 15036
rect 19740 14242 19796 14252
rect 20188 14868 20244 14878
rect 20188 14530 20244 14812
rect 20188 14478 20190 14530
rect 20242 14478 20244 14530
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19740 13860 19796 13870
rect 19740 12850 19796 13804
rect 20076 13524 20132 13534
rect 20076 13430 20132 13468
rect 20188 13076 20244 14478
rect 20188 13010 20244 13020
rect 19740 12798 19742 12850
rect 19794 12798 19796 12850
rect 19740 12786 19796 12798
rect 20188 12850 20244 12862
rect 20188 12798 20190 12850
rect 20242 12798 20244 12850
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19628 12348 20020 12404
rect 19628 12178 19684 12190
rect 19628 12126 19630 12178
rect 19682 12126 19684 12178
rect 19516 11394 19572 11406
rect 19516 11342 19518 11394
rect 19570 11342 19572 11394
rect 19516 11284 19572 11342
rect 19516 11218 19572 11228
rect 19404 10658 19460 10668
rect 19516 10612 19572 10622
rect 19516 10518 19572 10556
rect 19628 10164 19684 12126
rect 19852 11282 19908 11294
rect 19852 11230 19854 11282
rect 19906 11230 19908 11282
rect 19852 11172 19908 11230
rect 19964 11282 20020 12348
rect 20188 11956 20244 12798
rect 20300 12738 20356 15262
rect 20524 13858 20580 15596
rect 20748 15092 20804 22204
rect 20972 20020 21028 22540
rect 21196 22484 21252 24558
rect 21308 23716 21364 23726
rect 21308 23622 21364 23660
rect 21420 23380 21476 24780
rect 21868 24722 21924 24734
rect 21868 24670 21870 24722
rect 21922 24670 21924 24722
rect 21196 22418 21252 22428
rect 21308 23324 21476 23380
rect 21532 24612 21588 24622
rect 21532 24052 21588 24556
rect 21868 24612 21924 24670
rect 21868 24546 21924 24556
rect 21084 21700 21140 21710
rect 21084 21586 21140 21644
rect 21196 21700 21252 21710
rect 21308 21700 21364 23324
rect 21420 23156 21476 23166
rect 21420 23062 21476 23100
rect 21420 22372 21476 22382
rect 21420 22278 21476 22316
rect 21196 21698 21364 21700
rect 21196 21646 21198 21698
rect 21250 21646 21364 21698
rect 21196 21644 21364 21646
rect 21196 21634 21252 21644
rect 21084 21534 21086 21586
rect 21138 21534 21140 21586
rect 21084 21140 21140 21534
rect 21084 21074 21140 21084
rect 21084 20020 21140 20030
rect 20972 20018 21140 20020
rect 20972 19966 21086 20018
rect 21138 19966 21140 20018
rect 20972 19964 21140 19966
rect 20860 19908 20916 19918
rect 20860 19814 20916 19852
rect 20860 16884 20916 16894
rect 20860 16790 20916 16828
rect 20972 15148 21028 19964
rect 21084 19954 21140 19964
rect 21308 20018 21364 21644
rect 21308 19966 21310 20018
rect 21362 19966 21364 20018
rect 21308 19954 21364 19966
rect 21532 21364 21588 23996
rect 21756 24388 21812 24398
rect 21644 22370 21700 22382
rect 21644 22318 21646 22370
rect 21698 22318 21700 22370
rect 21644 22148 21700 22318
rect 21644 22082 21700 22092
rect 21420 19796 21476 19806
rect 21420 19346 21476 19740
rect 21420 19294 21422 19346
rect 21474 19294 21476 19346
rect 21420 19282 21476 19294
rect 21308 18452 21364 18462
rect 21308 18358 21364 18396
rect 21532 18228 21588 21308
rect 21644 20578 21700 20590
rect 21644 20526 21646 20578
rect 21698 20526 21700 20578
rect 21644 20468 21700 20526
rect 21644 20402 21700 20412
rect 21308 18172 21588 18228
rect 21196 17442 21252 17454
rect 21196 17390 21198 17442
rect 21250 17390 21252 17442
rect 21196 16996 21252 17390
rect 21308 17332 21364 18172
rect 21420 17556 21476 17566
rect 21420 17462 21476 17500
rect 21532 17556 21588 17566
rect 21532 17554 21700 17556
rect 21532 17502 21534 17554
rect 21586 17502 21700 17554
rect 21532 17500 21700 17502
rect 21532 17490 21588 17500
rect 21532 17332 21588 17342
rect 21308 17276 21476 17332
rect 21196 16930 21252 16940
rect 21308 16098 21364 16110
rect 21308 16046 21310 16098
rect 21362 16046 21364 16098
rect 21308 15540 21364 16046
rect 21420 15652 21476 17276
rect 21420 15586 21476 15596
rect 21308 15474 21364 15484
rect 21420 15428 21476 15438
rect 21420 15334 21476 15372
rect 20748 15026 20804 15036
rect 20860 15092 21028 15148
rect 21532 15148 21588 17276
rect 21644 16324 21700 17500
rect 21644 16258 21700 16268
rect 21084 15092 21140 15102
rect 21532 15092 21700 15148
rect 20748 14868 20804 14878
rect 20636 14644 20692 14654
rect 20636 14550 20692 14588
rect 20524 13806 20526 13858
rect 20578 13806 20580 13858
rect 20524 13794 20580 13806
rect 20636 13972 20692 13982
rect 20300 12686 20302 12738
rect 20354 12686 20356 12738
rect 20300 12674 20356 12686
rect 20412 13746 20468 13758
rect 20412 13694 20414 13746
rect 20466 13694 20468 13746
rect 20412 12292 20468 13694
rect 20636 13748 20692 13916
rect 20636 13682 20692 13692
rect 20748 13300 20804 14812
rect 20188 11890 20244 11900
rect 20300 12236 20412 12292
rect 19964 11230 19966 11282
rect 20018 11230 20020 11282
rect 19964 11218 20020 11230
rect 19852 11106 19908 11116
rect 20188 11172 20244 11182
rect 20188 11078 20244 11116
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20300 10948 20356 12236
rect 20412 12226 20468 12236
rect 20524 13244 20804 13300
rect 19836 10938 20100 10948
rect 20188 10892 20356 10948
rect 20412 12066 20468 12078
rect 20412 12014 20414 12066
rect 20466 12014 20468 12066
rect 19740 10836 19796 10846
rect 19796 10780 19908 10836
rect 19740 10770 19796 10780
rect 19628 10108 19796 10164
rect 19292 10098 19348 10108
rect 19292 9938 19348 9950
rect 19292 9886 19294 9938
rect 19346 9886 19348 9938
rect 19180 9826 19236 9838
rect 19180 9774 19182 9826
rect 19234 9774 19236 9826
rect 18844 9716 18900 9726
rect 18844 9714 19124 9716
rect 18844 9662 18846 9714
rect 18898 9662 19124 9714
rect 18844 9660 19124 9662
rect 18844 9650 18900 9660
rect 18732 9314 18788 9324
rect 18844 9492 18900 9502
rect 18732 9042 18788 9054
rect 18732 8990 18734 9042
rect 18786 8990 18788 9042
rect 18732 8484 18788 8990
rect 18732 8418 18788 8428
rect 18844 8146 18900 9436
rect 18956 9268 19012 9278
rect 19068 9268 19124 9660
rect 19180 9604 19236 9774
rect 19292 9828 19348 9886
rect 19292 9762 19348 9772
rect 19628 9716 19684 9726
rect 19628 9622 19684 9660
rect 19180 9538 19236 9548
rect 19404 9604 19460 9614
rect 19404 9510 19460 9548
rect 19740 9604 19796 10108
rect 19852 9604 19908 10780
rect 19964 10498 20020 10510
rect 19964 10446 19966 10498
rect 20018 10446 20020 10498
rect 19964 9940 20020 10446
rect 19964 9874 20020 9884
rect 20188 9826 20244 10892
rect 20300 10498 20356 10510
rect 20300 10446 20302 10498
rect 20354 10446 20356 10498
rect 20300 10164 20356 10446
rect 20300 10098 20356 10108
rect 20188 9774 20190 9826
rect 20242 9774 20244 9826
rect 20188 9762 20244 9774
rect 19964 9604 20020 9614
rect 19852 9548 19964 9604
rect 19740 9538 19796 9548
rect 19964 9538 20020 9548
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19068 9212 19460 9268
rect 18956 9174 19012 9212
rect 19404 9156 19460 9212
rect 19404 9154 20132 9156
rect 19404 9102 19406 9154
rect 19458 9102 20132 9154
rect 19404 9100 20132 9102
rect 19404 9090 19460 9100
rect 19068 9044 19124 9054
rect 19068 8950 19124 8988
rect 19292 9042 19348 9054
rect 19292 8990 19294 9042
rect 19346 8990 19348 9042
rect 19292 8932 19348 8990
rect 19404 8932 19460 8942
rect 19292 8876 19404 8932
rect 19404 8866 19460 8876
rect 18844 8094 18846 8146
rect 18898 8094 18900 8146
rect 18844 8082 18900 8094
rect 19180 8484 19236 8494
rect 18620 7644 18788 7700
rect 18620 7476 18676 7486
rect 18620 7382 18676 7420
rect 18508 7364 18564 7374
rect 18508 7270 18564 7308
rect 18396 6598 18452 6636
rect 18732 7252 18788 7644
rect 18732 6580 18788 7196
rect 18732 6514 18788 6524
rect 19068 6580 19124 6590
rect 18284 5854 18286 5906
rect 18338 5854 18340 5906
rect 18284 5348 18340 5854
rect 18508 6468 18564 6478
rect 18508 5908 18564 6412
rect 18620 6132 18676 6142
rect 18956 6132 19012 6142
rect 18620 6130 18788 6132
rect 18620 6078 18622 6130
rect 18674 6078 18788 6130
rect 18620 6076 18788 6078
rect 18620 6066 18676 6076
rect 18508 5814 18564 5852
rect 18284 5282 18340 5292
rect 18396 5236 18452 5246
rect 18396 5122 18452 5180
rect 18396 5070 18398 5122
rect 18450 5070 18452 5122
rect 18396 5058 18452 5070
rect 18620 5124 18676 5134
rect 18620 5030 18676 5068
rect 18732 5012 18788 6076
rect 18956 6038 19012 6076
rect 18956 5124 19012 5134
rect 19068 5124 19124 6524
rect 18956 5122 19124 5124
rect 18956 5070 18958 5122
rect 19010 5070 19124 5122
rect 18956 5068 19124 5070
rect 18956 5058 19012 5068
rect 18732 4946 18788 4956
rect 19180 5010 19236 8428
rect 19628 8484 19684 8494
rect 19628 7700 19684 8428
rect 20076 8258 20132 9100
rect 20076 8206 20078 8258
rect 20130 8206 20132 8258
rect 20076 8194 20132 8206
rect 20188 8820 20244 8830
rect 20188 8484 20244 8764
rect 19964 8148 20020 8158
rect 19964 8054 20020 8092
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19852 7700 19908 7710
rect 19628 7698 19908 7700
rect 19628 7646 19854 7698
rect 19906 7646 19908 7698
rect 19628 7644 19908 7646
rect 19852 7634 19908 7644
rect 20076 7700 20132 7710
rect 20076 7606 20132 7644
rect 19964 7588 20020 7598
rect 19292 7532 19796 7588
rect 19292 7474 19348 7532
rect 19292 7422 19294 7474
rect 19346 7422 19348 7474
rect 19292 7410 19348 7422
rect 19740 7476 19796 7532
rect 19964 7476 20020 7532
rect 20188 7586 20244 8428
rect 20412 7700 20468 12014
rect 20524 10612 20580 13244
rect 20860 13188 20916 15092
rect 21084 14420 21140 15036
rect 21084 13970 21140 14364
rect 21084 13918 21086 13970
rect 21138 13918 21140 13970
rect 21084 13906 21140 13918
rect 21196 14532 21252 14542
rect 20972 13748 21028 13758
rect 20972 13654 21028 13692
rect 20636 13132 20916 13188
rect 20636 10836 20692 13132
rect 20748 12964 20804 12974
rect 20748 11732 20804 12908
rect 20860 11844 20916 11854
rect 20916 11788 21028 11844
rect 20860 11778 20916 11788
rect 20748 11506 20804 11676
rect 20748 11454 20750 11506
rect 20802 11454 20804 11506
rect 20748 11442 20804 11454
rect 20636 10780 20916 10836
rect 20524 10546 20580 10556
rect 20748 10610 20804 10622
rect 20748 10558 20750 10610
rect 20802 10558 20804 10610
rect 20748 10052 20804 10558
rect 20748 9986 20804 9996
rect 20636 9828 20692 9838
rect 20636 9734 20692 9772
rect 20412 7634 20468 7644
rect 20524 9716 20580 9726
rect 20524 9602 20580 9660
rect 20524 9550 20526 9602
rect 20578 9550 20580 9602
rect 20524 8932 20580 9550
rect 20748 9604 20804 9614
rect 20748 9510 20804 9548
rect 20188 7534 20190 7586
rect 20242 7534 20244 7586
rect 20188 7522 20244 7534
rect 19740 7420 20020 7476
rect 20300 7476 20356 7486
rect 20524 7476 20580 8876
rect 19404 7364 19460 7374
rect 19404 7270 19460 7308
rect 19292 7252 19348 7262
rect 19292 6690 19348 7196
rect 19292 6638 19294 6690
rect 19346 6638 19348 6690
rect 19292 6626 19348 6638
rect 19628 7028 19684 7038
rect 19628 6690 19684 6972
rect 19964 6804 20020 6814
rect 19964 6802 20244 6804
rect 19964 6750 19966 6802
rect 20018 6750 20244 6802
rect 19964 6748 20244 6750
rect 19964 6738 20020 6748
rect 19628 6638 19630 6690
rect 19682 6638 19684 6690
rect 19516 5908 19572 5918
rect 19516 5814 19572 5852
rect 19628 5460 19684 6638
rect 20188 6690 20244 6748
rect 20188 6638 20190 6690
rect 20242 6638 20244 6690
rect 20188 6626 20244 6638
rect 19852 6580 19908 6590
rect 19852 6486 19908 6524
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 20188 6132 20244 6142
rect 20188 6038 20244 6076
rect 19852 6020 19908 6030
rect 19852 5926 19908 5964
rect 20300 5908 20356 7420
rect 20076 5852 20356 5908
rect 20412 7420 20580 7476
rect 20636 7700 20692 7710
rect 20860 7700 20916 10780
rect 20972 7812 21028 11788
rect 21084 11172 21140 11182
rect 21084 10610 21140 11116
rect 21084 10558 21086 10610
rect 21138 10558 21140 10610
rect 21084 10388 21140 10558
rect 21084 10322 21140 10332
rect 21196 10052 21252 14476
rect 21532 14532 21588 14542
rect 21532 14438 21588 14476
rect 21308 14196 21364 14206
rect 21308 13970 21364 14140
rect 21308 13918 21310 13970
rect 21362 13918 21364 13970
rect 21308 13906 21364 13918
rect 21532 13972 21588 13982
rect 21532 13858 21588 13916
rect 21532 13806 21534 13858
rect 21586 13806 21588 13858
rect 21532 13794 21588 13806
rect 21308 12180 21364 12190
rect 21644 12180 21700 15092
rect 21756 14868 21812 24332
rect 22092 24164 22148 24174
rect 22092 23938 22148 24108
rect 22092 23886 22094 23938
rect 22146 23886 22148 23938
rect 22092 23874 22148 23886
rect 21868 23604 21924 23614
rect 21868 23378 21924 23548
rect 21868 23326 21870 23378
rect 21922 23326 21924 23378
rect 21868 23314 21924 23326
rect 22316 22372 22372 24892
rect 22428 24722 22484 27132
rect 22428 24670 22430 24722
rect 22482 24670 22484 24722
rect 22428 24658 22484 24670
rect 22540 25284 22596 25294
rect 22540 23938 22596 25228
rect 22540 23886 22542 23938
rect 22594 23886 22596 23938
rect 22540 23874 22596 23886
rect 22428 23380 22484 23390
rect 22428 23266 22484 23324
rect 22428 23214 22430 23266
rect 22482 23214 22484 23266
rect 22428 23202 22484 23214
rect 22652 23266 22708 28588
rect 22764 28550 22820 28588
rect 23100 28420 23156 28430
rect 22764 28084 22820 28094
rect 22764 27188 22820 28028
rect 22764 27094 22820 27132
rect 22988 26516 23044 26526
rect 22988 26290 23044 26460
rect 22988 26238 22990 26290
rect 23042 26238 23044 26290
rect 22988 26226 23044 26238
rect 22764 25620 22820 25630
rect 22764 25618 22932 25620
rect 22764 25566 22766 25618
rect 22818 25566 22932 25618
rect 22764 25564 22932 25566
rect 22764 25554 22820 25564
rect 22652 23214 22654 23266
rect 22706 23214 22708 23266
rect 22316 22306 22372 22316
rect 22428 21810 22484 21822
rect 22428 21758 22430 21810
rect 22482 21758 22484 21810
rect 21868 21586 21924 21598
rect 21868 21534 21870 21586
rect 21922 21534 21924 21586
rect 21868 21476 21924 21534
rect 22428 21588 22484 21758
rect 22428 21522 22484 21532
rect 21868 21410 21924 21420
rect 22204 20804 22260 20814
rect 22092 20802 22260 20804
rect 22092 20750 22206 20802
rect 22258 20750 22260 20802
rect 22092 20748 22260 20750
rect 22092 20242 22148 20748
rect 22204 20738 22260 20748
rect 22316 20690 22372 20702
rect 22316 20638 22318 20690
rect 22370 20638 22372 20690
rect 22316 20244 22372 20638
rect 22428 20578 22484 20590
rect 22428 20526 22430 20578
rect 22482 20526 22484 20578
rect 22428 20356 22484 20526
rect 22428 20290 22484 20300
rect 22540 20580 22596 20590
rect 22092 20190 22094 20242
rect 22146 20190 22148 20242
rect 22092 20178 22148 20190
rect 22204 20188 22372 20244
rect 21868 19234 21924 19246
rect 21868 19182 21870 19234
rect 21922 19182 21924 19234
rect 21868 18676 21924 19182
rect 21868 18610 21924 18620
rect 22204 17892 22260 20188
rect 22428 20132 22484 20142
rect 22428 20038 22484 20076
rect 22316 20018 22372 20030
rect 22316 19966 22318 20018
rect 22370 19966 22372 20018
rect 22316 19348 22372 19966
rect 22316 19282 22372 19292
rect 22316 19124 22372 19134
rect 22316 19030 22372 19068
rect 22540 18900 22596 20524
rect 22652 20468 22708 23214
rect 22876 23268 22932 25564
rect 23100 24724 23156 28364
rect 24556 28084 24612 28590
rect 24668 28532 24724 28542
rect 24668 28438 24724 28476
rect 24668 28084 24724 28094
rect 24556 28028 24668 28084
rect 24668 27990 24724 28028
rect 23548 27858 23604 27870
rect 23548 27806 23550 27858
rect 23602 27806 23604 27858
rect 23548 27524 23604 27806
rect 23212 27074 23268 27086
rect 23212 27022 23214 27074
rect 23266 27022 23268 27074
rect 23212 25508 23268 27022
rect 23212 25414 23268 25452
rect 23324 26964 23380 26974
rect 23212 24948 23268 24958
rect 23324 24948 23380 26908
rect 23548 26962 23604 27468
rect 23548 26910 23550 26962
rect 23602 26910 23604 26962
rect 23548 26898 23604 26910
rect 23996 27746 24052 27758
rect 23996 27694 23998 27746
rect 24050 27694 24052 27746
rect 23772 26178 23828 26190
rect 23772 26126 23774 26178
rect 23826 26126 23828 26178
rect 23268 24892 23380 24948
rect 23436 25956 23492 25966
rect 23212 24882 23268 24892
rect 23436 24834 23492 25900
rect 23436 24782 23438 24834
rect 23490 24782 23492 24834
rect 23436 24770 23492 24782
rect 23212 24724 23268 24734
rect 23100 24722 23268 24724
rect 23100 24670 23214 24722
rect 23266 24670 23268 24722
rect 23100 24668 23268 24670
rect 23212 24500 23268 24668
rect 23324 24612 23380 24622
rect 23324 24518 23380 24556
rect 22988 23938 23044 23950
rect 22988 23886 22990 23938
rect 23042 23886 23044 23938
rect 22988 23492 23044 23886
rect 22988 23426 23044 23436
rect 22876 23212 23156 23268
rect 22764 23044 22820 23054
rect 22764 22950 22820 22988
rect 22764 20468 22820 20478
rect 22652 20412 22764 20468
rect 22764 20402 22820 20412
rect 22876 19908 22932 23212
rect 23100 23154 23156 23212
rect 23100 23102 23102 23154
rect 23154 23102 23156 23154
rect 23100 23090 23156 23102
rect 22988 22596 23044 22606
rect 22988 22260 23044 22540
rect 22988 20804 23044 22204
rect 23100 21588 23156 21598
rect 23100 21494 23156 21532
rect 22988 20748 23156 20804
rect 22540 18834 22596 18844
rect 22764 19852 22932 19908
rect 22764 19234 22820 19852
rect 22988 19460 23044 19470
rect 22764 19182 22766 19234
rect 22818 19182 22820 19234
rect 22428 18452 22484 18462
rect 22652 18452 22708 18462
rect 22428 18358 22484 18396
rect 22540 18450 22708 18452
rect 22540 18398 22654 18450
rect 22706 18398 22708 18450
rect 22540 18396 22708 18398
rect 21868 17836 22260 17892
rect 22540 18228 22596 18396
rect 22652 18386 22708 18396
rect 21868 16548 21924 17836
rect 21868 16482 21924 16492
rect 21980 17668 22036 17678
rect 21980 15988 22036 17612
rect 21980 15922 22036 15932
rect 22092 17666 22148 17678
rect 22092 17614 22094 17666
rect 22146 17614 22148 17666
rect 22092 15876 22148 17614
rect 22540 17554 22596 18172
rect 22540 17502 22542 17554
rect 22594 17502 22596 17554
rect 22540 17490 22596 17502
rect 22764 16884 22820 19182
rect 22092 15810 22148 15820
rect 22204 16882 22820 16884
rect 22204 16830 22766 16882
rect 22818 16830 22820 16882
rect 22204 16828 22820 16830
rect 21980 15764 22036 15774
rect 21756 14802 21812 14812
rect 21868 15314 21924 15326
rect 21868 15262 21870 15314
rect 21922 15262 21924 15314
rect 21868 14754 21924 15262
rect 21868 14702 21870 14754
rect 21922 14702 21924 14754
rect 21868 14690 21924 14702
rect 21980 14642 22036 15708
rect 22204 15148 22260 16828
rect 22764 16818 22820 16828
rect 22876 19236 22932 19246
rect 22876 19122 22932 19180
rect 22988 19234 23044 19404
rect 22988 19182 22990 19234
rect 23042 19182 23044 19234
rect 22988 19170 23044 19182
rect 22876 19070 22878 19122
rect 22930 19070 22932 19122
rect 21980 14590 21982 14642
rect 22034 14590 22036 14642
rect 21868 13746 21924 13758
rect 21868 13694 21870 13746
rect 21922 13694 21924 13746
rect 21868 13636 21924 13694
rect 21868 13570 21924 13580
rect 21756 12964 21812 12974
rect 21756 12962 21924 12964
rect 21756 12910 21758 12962
rect 21810 12910 21924 12962
rect 21756 12908 21924 12910
rect 21756 12898 21812 12908
rect 21756 12180 21812 12190
rect 21644 12124 21756 12180
rect 21308 12086 21364 12124
rect 21756 12114 21812 12124
rect 21868 11844 21924 12908
rect 21980 12628 22036 14590
rect 21980 12562 22036 12572
rect 22092 15092 22260 15148
rect 22316 16212 22372 16222
rect 21980 12290 22036 12302
rect 21980 12238 21982 12290
rect 22034 12238 22036 12290
rect 21980 11956 22036 12238
rect 21980 11890 22036 11900
rect 21868 11778 21924 11788
rect 21756 11506 21812 11518
rect 21756 11454 21758 11506
rect 21810 11454 21812 11506
rect 21756 11060 21812 11454
rect 22092 11394 22148 15092
rect 22316 14420 22372 16156
rect 22428 16100 22484 16110
rect 22764 16100 22820 16110
rect 22428 16006 22484 16044
rect 22540 16044 22764 16100
rect 22540 15876 22596 16044
rect 22764 16034 22820 16044
rect 22092 11342 22094 11394
rect 22146 11342 22148 11394
rect 22092 11330 22148 11342
rect 22204 14084 22260 14094
rect 21532 11004 21756 11060
rect 21196 9996 21476 10052
rect 21308 9826 21364 9838
rect 21308 9774 21310 9826
rect 21362 9774 21364 9826
rect 21084 9716 21140 9726
rect 21084 8596 21140 9660
rect 21084 8530 21140 8540
rect 20972 7746 21028 7756
rect 20636 7474 20692 7644
rect 20636 7422 20638 7474
rect 20690 7422 20692 7474
rect 20412 6578 20468 7420
rect 20636 7410 20692 7422
rect 20748 7644 20916 7700
rect 20748 7476 20804 7644
rect 20860 7476 20916 7486
rect 20748 7474 20916 7476
rect 20748 7422 20862 7474
rect 20914 7422 20916 7474
rect 20748 7420 20916 7422
rect 20748 6804 20804 7420
rect 20860 7410 20916 7420
rect 21084 7250 21140 7262
rect 21084 7198 21086 7250
rect 21138 7198 21140 7250
rect 20748 6738 20804 6748
rect 20860 6916 20916 6926
rect 20412 6526 20414 6578
rect 20466 6526 20468 6578
rect 20412 5908 20468 6526
rect 20524 6692 20580 6702
rect 20524 6244 20580 6636
rect 20748 6578 20804 6590
rect 20748 6526 20750 6578
rect 20802 6526 20804 6578
rect 20636 6468 20692 6478
rect 20636 6374 20692 6412
rect 20524 6188 20692 6244
rect 20636 6018 20692 6188
rect 20636 5966 20638 6018
rect 20690 5966 20692 6018
rect 20636 5954 20692 5966
rect 19180 4958 19182 5010
rect 19234 4958 19236 5010
rect 19068 4898 19124 4910
rect 19068 4846 19070 4898
rect 19122 4846 19124 4898
rect 18396 4564 18452 4574
rect 18396 4470 18452 4508
rect 18284 4452 18340 4462
rect 18172 4396 18284 4452
rect 18284 4386 18340 4396
rect 18844 4452 18900 4462
rect 18844 4358 18900 4396
rect 19068 4450 19124 4846
rect 19180 4676 19236 4958
rect 19292 5404 19684 5460
rect 19852 5684 19908 5694
rect 19292 4900 19348 5404
rect 19740 5348 19796 5358
rect 19628 5292 19740 5348
rect 19516 5236 19572 5246
rect 19292 4834 19348 4844
rect 19404 5180 19516 5236
rect 19180 4610 19236 4620
rect 19068 4398 19070 4450
rect 19122 4398 19124 4450
rect 19068 4386 19124 4398
rect 19292 4452 19348 4462
rect 18620 4340 18676 4350
rect 17724 3614 17726 3666
rect 17778 3614 17780 3666
rect 17724 3602 17780 3614
rect 18172 3778 18228 3790
rect 18172 3726 18174 3778
rect 18226 3726 18228 3778
rect 18172 3666 18228 3726
rect 18172 3614 18174 3666
rect 18226 3614 18228 3666
rect 18172 3602 18228 3614
rect 18620 3666 18676 4284
rect 19292 3892 19348 4396
rect 19404 4228 19460 5180
rect 19516 5170 19572 5180
rect 19516 5010 19572 5022
rect 19516 4958 19518 5010
rect 19570 4958 19572 5010
rect 19516 4900 19572 4958
rect 19516 4834 19572 4844
rect 19628 4452 19684 5292
rect 19740 5282 19796 5292
rect 19852 5346 19908 5628
rect 19852 5294 19854 5346
rect 19906 5294 19908 5346
rect 19852 5282 19908 5294
rect 20076 5236 20132 5852
rect 20412 5842 20468 5852
rect 20524 5906 20580 5918
rect 20524 5854 20526 5906
rect 20578 5854 20580 5906
rect 20524 5796 20580 5854
rect 20524 5730 20580 5740
rect 19740 5122 19796 5134
rect 19740 5070 19742 5122
rect 19794 5070 19796 5122
rect 19740 4900 19796 5070
rect 20076 4900 20132 5180
rect 20300 5572 20356 5582
rect 19740 4844 20132 4900
rect 20188 4900 20244 4910
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19964 4564 20020 4574
rect 19964 4470 20020 4508
rect 19628 4396 19796 4452
rect 19628 4228 19684 4238
rect 19404 4226 19684 4228
rect 19404 4174 19630 4226
rect 19682 4174 19684 4226
rect 19404 4172 19684 4174
rect 19628 4162 19684 4172
rect 19292 3826 19348 3836
rect 18620 3614 18622 3666
rect 18674 3614 18676 3666
rect 18620 3602 18676 3614
rect 19180 3668 19236 3678
rect 19236 3612 19348 3668
rect 19180 3602 19236 3612
rect 19292 3554 19348 3612
rect 19292 3502 19294 3554
rect 19346 3502 19348 3554
rect 19292 3490 19348 3502
rect 19740 3666 19796 4396
rect 19852 4340 19908 4350
rect 20188 4340 20244 4844
rect 19852 4338 20244 4340
rect 19852 4286 19854 4338
rect 19906 4286 20244 4338
rect 19852 4284 20244 4286
rect 19852 4274 19908 4284
rect 19740 3614 19742 3666
rect 19794 3614 19796 3666
rect 19740 3332 19796 3614
rect 20188 3668 20244 3678
rect 20300 3668 20356 5516
rect 20524 5460 20580 5470
rect 20524 5346 20580 5404
rect 20524 5294 20526 5346
rect 20578 5294 20580 5346
rect 20524 5282 20580 5294
rect 20748 5348 20804 6526
rect 20860 5684 20916 6860
rect 20860 5618 20916 5628
rect 21084 6356 21140 7198
rect 21084 5572 21140 6300
rect 21084 5506 21140 5516
rect 21196 6804 21252 6814
rect 20748 5282 20804 5292
rect 20636 5236 20692 5246
rect 20636 5012 20692 5180
rect 20748 5012 20804 5022
rect 21196 5012 21252 6748
rect 21308 6132 21364 9774
rect 21420 8372 21476 9996
rect 21532 8372 21588 11004
rect 21756 10994 21812 11004
rect 22204 10610 22260 14028
rect 22204 10558 22206 10610
rect 22258 10558 22260 10610
rect 22204 10546 22260 10558
rect 21980 10498 22036 10510
rect 21980 10446 21982 10498
rect 22034 10446 22036 10498
rect 21644 10052 21700 10062
rect 21644 9826 21700 9996
rect 21756 9940 21812 9950
rect 21756 9846 21812 9884
rect 21644 9774 21646 9826
rect 21698 9774 21700 9826
rect 21644 9762 21700 9774
rect 21868 9828 21924 9838
rect 21980 9828 22036 10446
rect 21868 9826 22036 9828
rect 21868 9774 21870 9826
rect 21922 9774 22036 9826
rect 21868 9772 22036 9774
rect 21868 9762 21924 9772
rect 21980 9604 22036 9772
rect 21980 9538 22036 9548
rect 22092 10164 22148 10174
rect 21644 9042 21700 9054
rect 21644 8990 21646 9042
rect 21698 8990 21700 9042
rect 21644 8932 21700 8990
rect 21644 8866 21700 8876
rect 21980 9042 22036 9054
rect 21980 8990 21982 9042
rect 22034 8990 22036 9042
rect 21980 8484 22036 8990
rect 21980 8418 22036 8428
rect 21532 8316 21924 8372
rect 21420 8278 21476 8316
rect 21532 8148 21588 8158
rect 21532 7698 21588 8092
rect 21532 7646 21534 7698
rect 21586 7646 21588 7698
rect 21532 7634 21588 7646
rect 21868 7700 21924 8316
rect 21868 7606 21924 7644
rect 21644 7476 21700 7486
rect 21644 7382 21700 7420
rect 21980 7474 22036 7486
rect 21980 7422 21982 7474
rect 22034 7422 22036 7474
rect 21980 7252 22036 7422
rect 21980 7186 22036 7196
rect 21756 7028 21812 7038
rect 21420 6692 21476 6702
rect 21420 6598 21476 6636
rect 21644 6580 21700 6590
rect 21532 6132 21588 6142
rect 21308 6130 21588 6132
rect 21308 6078 21534 6130
rect 21586 6078 21588 6130
rect 21308 6076 21588 6078
rect 21532 5796 21588 6076
rect 21644 5908 21700 6524
rect 21644 5814 21700 5852
rect 21532 5730 21588 5740
rect 20636 5010 20804 5012
rect 20636 4958 20750 5010
rect 20802 4958 20804 5010
rect 20636 4956 20804 4958
rect 20524 4226 20580 4238
rect 20524 4174 20526 4226
rect 20578 4174 20580 4226
rect 20524 4116 20580 4174
rect 20524 4050 20580 4060
rect 20748 3778 20804 4956
rect 20748 3726 20750 3778
rect 20802 3726 20804 3778
rect 20748 3714 20804 3726
rect 20972 4956 21252 5012
rect 21308 5684 21364 5694
rect 20188 3666 20356 3668
rect 20188 3614 20190 3666
rect 20242 3614 20356 3666
rect 20188 3612 20356 3614
rect 20972 3666 21028 4956
rect 21084 4564 21140 4574
rect 21308 4564 21364 5628
rect 21756 5122 21812 6972
rect 22092 6916 22148 10108
rect 22204 9826 22260 9838
rect 22204 9774 22206 9826
rect 22258 9774 22260 9826
rect 22204 7028 22260 9774
rect 22316 8484 22372 14364
rect 22428 15820 22596 15876
rect 22428 13860 22484 15820
rect 22540 15652 22596 15662
rect 22540 14756 22596 15596
rect 22764 15428 22820 15466
rect 22764 15362 22820 15372
rect 22652 15314 22708 15326
rect 22652 15262 22654 15314
rect 22706 15262 22708 15314
rect 22652 14980 22708 15262
rect 22764 15204 22820 15242
rect 22764 15138 22820 15148
rect 22652 14914 22708 14924
rect 22764 14756 22820 14766
rect 22540 14700 22708 14756
rect 22428 13794 22484 13804
rect 22428 12964 22484 12974
rect 22428 12870 22484 12908
rect 22540 12404 22596 12414
rect 22652 12404 22708 14700
rect 22764 14530 22820 14700
rect 22764 14478 22766 14530
rect 22818 14478 22820 14530
rect 22764 14466 22820 14478
rect 22876 14420 22932 19070
rect 22988 18452 23044 18462
rect 22988 17556 23044 18396
rect 23100 17666 23156 20748
rect 23212 17892 23268 24444
rect 23772 24164 23828 26126
rect 23996 26068 24052 27694
rect 23996 26002 24052 26012
rect 24220 27186 24276 27198
rect 24220 27134 24222 27186
rect 24274 27134 24276 27186
rect 23884 25508 23940 25518
rect 23940 25452 24164 25508
rect 23884 25414 23940 25452
rect 24108 24834 24164 25452
rect 24108 24782 24110 24834
rect 24162 24782 24164 24834
rect 24108 24770 24164 24782
rect 23772 24098 23828 24108
rect 23996 23940 24052 23950
rect 24220 23940 24276 27134
rect 24780 26908 24836 29150
rect 25228 28756 25284 28766
rect 25228 28754 25620 28756
rect 25228 28702 25230 28754
rect 25282 28702 25620 28754
rect 25228 28700 25620 28702
rect 25228 28690 25284 28700
rect 25564 28644 25620 28700
rect 26124 28644 26180 28654
rect 25564 28642 25956 28644
rect 25564 28590 25566 28642
rect 25618 28590 25956 28642
rect 25564 28588 25956 28590
rect 25564 28578 25620 28588
rect 25676 28084 25732 28094
rect 25676 27858 25732 28028
rect 25676 27806 25678 27858
rect 25730 27806 25732 27858
rect 25676 27794 25732 27806
rect 25340 27746 25396 27758
rect 25340 27694 25342 27746
rect 25394 27694 25396 27746
rect 24332 26852 24388 26862
rect 24780 26852 25060 26908
rect 24332 26402 24388 26796
rect 24332 26350 24334 26402
rect 24386 26350 24388 26402
rect 24332 26338 24388 26350
rect 24780 26404 24836 26414
rect 24444 26292 24500 26302
rect 24444 26290 24724 26292
rect 24444 26238 24446 26290
rect 24498 26238 24724 26290
rect 24444 26236 24724 26238
rect 24444 26226 24500 26236
rect 24332 26180 24388 26190
rect 24332 25284 24388 26124
rect 24556 25284 24612 25294
rect 24332 25282 24612 25284
rect 24332 25230 24558 25282
rect 24610 25230 24612 25282
rect 24332 25228 24612 25230
rect 24444 23940 24500 23950
rect 24220 23938 24500 23940
rect 24220 23886 24446 23938
rect 24498 23886 24500 23938
rect 24220 23884 24500 23886
rect 23996 23826 24052 23884
rect 23996 23774 23998 23826
rect 24050 23774 24052 23826
rect 23996 23762 24052 23774
rect 23436 23492 23492 23502
rect 23324 22930 23380 22942
rect 23324 22878 23326 22930
rect 23378 22878 23380 22930
rect 23324 22708 23380 22878
rect 23324 22642 23380 22652
rect 23436 22372 23492 23436
rect 24444 23492 24500 23884
rect 24444 23426 24500 23436
rect 24332 23154 24388 23166
rect 24332 23102 24334 23154
rect 24386 23102 24388 23154
rect 23660 22932 23716 22942
rect 23660 22930 23828 22932
rect 23660 22878 23662 22930
rect 23714 22878 23828 22930
rect 23660 22876 23828 22878
rect 23660 22866 23716 22876
rect 23436 22306 23492 22316
rect 23548 22370 23604 22382
rect 23548 22318 23550 22370
rect 23602 22318 23604 22370
rect 23548 21700 23604 22318
rect 23604 21644 23716 21700
rect 23548 21634 23604 21644
rect 23436 21588 23492 21598
rect 23436 21494 23492 21532
rect 23660 21028 23716 21644
rect 23772 21252 23828 22876
rect 24332 21812 24388 23102
rect 24332 21746 24388 21756
rect 24444 23042 24500 23054
rect 24444 22990 24446 23042
rect 24498 22990 24500 23042
rect 24332 21588 24388 21598
rect 24444 21588 24500 22990
rect 24332 21586 24500 21588
rect 24332 21534 24334 21586
rect 24386 21534 24500 21586
rect 24332 21532 24500 21534
rect 23884 21476 23940 21486
rect 23884 21382 23940 21420
rect 24220 21364 24276 21374
rect 24220 21270 24276 21308
rect 23772 21196 24052 21252
rect 23660 20972 23940 21028
rect 23772 20804 23828 20814
rect 23324 20802 23828 20804
rect 23324 20750 23774 20802
rect 23826 20750 23828 20802
rect 23324 20748 23828 20750
rect 23324 20242 23380 20748
rect 23772 20738 23828 20748
rect 23324 20190 23326 20242
rect 23378 20190 23380 20242
rect 23324 20178 23380 20190
rect 23436 20020 23492 20030
rect 23436 19926 23492 19964
rect 23884 19458 23940 20972
rect 23996 20018 24052 21196
rect 24220 20132 24276 20142
rect 24220 20038 24276 20076
rect 23996 19966 23998 20018
rect 24050 19966 24052 20018
rect 23996 19954 24052 19966
rect 23884 19406 23886 19458
rect 23938 19406 23940 19458
rect 23884 19394 23940 19406
rect 23996 19572 24052 19582
rect 23996 19458 24052 19516
rect 23996 19406 23998 19458
rect 24050 19406 24052 19458
rect 23996 19394 24052 19406
rect 24220 19572 24276 19582
rect 24220 19458 24276 19516
rect 24220 19406 24222 19458
rect 24274 19406 24276 19458
rect 24220 19394 24276 19406
rect 23884 19124 23940 19134
rect 23436 19010 23492 19022
rect 23436 18958 23438 19010
rect 23490 18958 23492 19010
rect 23324 18900 23380 18910
rect 23324 18564 23380 18844
rect 23436 18676 23492 18958
rect 23884 19010 23940 19068
rect 23884 18958 23886 19010
rect 23938 18958 23940 19010
rect 23884 18946 23940 18958
rect 23436 18620 23604 18676
rect 23324 18508 23492 18564
rect 23324 18340 23380 18350
rect 23324 18246 23380 18284
rect 23324 17892 23380 17902
rect 23212 17836 23324 17892
rect 23324 17826 23380 17836
rect 23436 17668 23492 18508
rect 23100 17614 23102 17666
rect 23154 17614 23156 17666
rect 23100 17602 23156 17614
rect 23324 17612 23492 17668
rect 23548 17668 23604 18620
rect 24220 18674 24276 18686
rect 24220 18622 24222 18674
rect 24274 18622 24276 18674
rect 23772 18564 23828 18574
rect 23772 18452 23828 18508
rect 23772 18450 23940 18452
rect 23772 18398 23774 18450
rect 23826 18398 23940 18450
rect 23772 18396 23940 18398
rect 23772 18386 23828 18396
rect 23772 18228 23828 18238
rect 23772 18134 23828 18172
rect 23772 18004 23828 18014
rect 23772 17780 23828 17948
rect 23772 17686 23828 17724
rect 22988 17490 23044 17500
rect 23100 17442 23156 17454
rect 23100 17390 23102 17442
rect 23154 17390 23156 17442
rect 23100 16884 23156 17390
rect 23100 16818 23156 16828
rect 23324 16100 23380 17612
rect 23548 17602 23604 17612
rect 23772 16996 23828 17006
rect 23772 16902 23828 16940
rect 23436 16212 23492 16222
rect 23436 16118 23492 16156
rect 23324 16006 23380 16044
rect 23884 16100 23940 18396
rect 24220 17444 24276 18622
rect 24332 18452 24388 21532
rect 24556 20580 24612 25228
rect 24668 25284 24724 26236
rect 24668 24946 24724 25228
rect 24668 24894 24670 24946
rect 24722 24894 24724 24946
rect 24668 24882 24724 24894
rect 24668 23266 24724 23278
rect 24668 23214 24670 23266
rect 24722 23214 24724 23266
rect 24668 23156 24724 23214
rect 24668 23090 24724 23100
rect 24668 22260 24724 22270
rect 24780 22260 24836 26348
rect 24668 22258 24836 22260
rect 24668 22206 24670 22258
rect 24722 22206 24836 22258
rect 24668 22204 24836 22206
rect 24668 22194 24724 22204
rect 24892 22148 24948 22158
rect 24892 22054 24948 22092
rect 24556 20514 24612 20524
rect 24444 20018 24500 20030
rect 24444 19966 24446 20018
rect 24498 19966 24500 20018
rect 24444 18674 24500 19966
rect 24444 18622 24446 18674
rect 24498 18622 24500 18674
rect 24444 18610 24500 18622
rect 24556 20018 24612 20030
rect 24556 19966 24558 20018
rect 24610 19966 24612 20018
rect 24332 18396 24500 18452
rect 24332 17668 24388 17678
rect 24332 17574 24388 17612
rect 24220 17378 24276 17388
rect 24332 17108 24388 17118
rect 24444 17108 24500 18396
rect 24556 18340 24612 19966
rect 25004 19236 25060 26852
rect 25228 25844 25284 25854
rect 25116 25508 25172 25518
rect 25116 25414 25172 25452
rect 25228 24948 25284 25788
rect 25340 25284 25396 27694
rect 25340 25218 25396 25228
rect 25452 27524 25508 27534
rect 25452 27074 25508 27468
rect 25452 27022 25454 27074
rect 25506 27022 25508 27074
rect 25228 24882 25284 24892
rect 25340 24724 25396 24734
rect 25340 23492 25396 24668
rect 25452 23940 25508 27022
rect 25788 26964 25844 27002
rect 25788 26898 25844 26908
rect 25788 26068 25844 26078
rect 25564 24724 25620 24734
rect 25564 24630 25620 24668
rect 25788 24052 25844 26012
rect 25900 25618 25956 28588
rect 26124 28550 26180 28588
rect 26124 28084 26180 28094
rect 26124 27970 26180 28028
rect 26908 28084 26964 28094
rect 27692 28084 27748 28094
rect 26908 27990 26964 28028
rect 27580 28028 27692 28084
rect 26124 27918 26126 27970
rect 26178 27918 26180 27970
rect 26124 27906 26180 27918
rect 27468 27860 27524 27870
rect 26460 27746 26516 27758
rect 26460 27694 26462 27746
rect 26514 27694 26516 27746
rect 26236 27188 26292 27198
rect 26236 26908 26292 27132
rect 26460 27076 26516 27694
rect 26460 27010 26516 27020
rect 27132 27076 27188 27086
rect 27132 26962 27188 27020
rect 27132 26910 27134 26962
rect 27186 26910 27188 26962
rect 26236 26852 26516 26908
rect 27132 26898 27188 26910
rect 27244 27074 27300 27086
rect 27244 27022 27246 27074
rect 27298 27022 27300 27074
rect 26460 26290 26516 26852
rect 27244 26852 27300 27022
rect 27244 26786 27300 26796
rect 26460 26238 26462 26290
rect 26514 26238 26516 26290
rect 26460 26226 26516 26238
rect 26348 26180 26404 26190
rect 25900 25566 25902 25618
rect 25954 25566 25956 25618
rect 25900 25554 25956 25566
rect 26012 26178 26404 26180
rect 26012 26126 26350 26178
rect 26402 26126 26404 26178
rect 26012 26124 26404 26126
rect 26012 25956 26068 26124
rect 26348 26114 26404 26124
rect 26012 24610 26068 25900
rect 27356 26068 27412 26078
rect 26124 25506 26180 25518
rect 26124 25454 26126 25506
rect 26178 25454 26180 25506
rect 26124 25396 26180 25454
rect 26124 25330 26180 25340
rect 26012 24558 26014 24610
rect 26066 24558 26068 24610
rect 26012 24546 26068 24558
rect 26572 24722 26628 24734
rect 26572 24670 26574 24722
rect 26626 24670 26628 24722
rect 26572 24612 26628 24670
rect 26460 24498 26516 24510
rect 26460 24446 26462 24498
rect 26514 24446 26516 24498
rect 25788 23996 25956 24052
rect 25452 23884 25844 23940
rect 25452 23716 25508 23726
rect 25452 23622 25508 23660
rect 25564 23492 25620 23502
rect 25340 23436 25508 23492
rect 25340 23044 25396 23054
rect 25340 22950 25396 22988
rect 25452 22482 25508 23436
rect 25452 22430 25454 22482
rect 25506 22430 25508 22482
rect 25452 22418 25508 22430
rect 25228 21586 25284 21598
rect 25228 21534 25230 21586
rect 25282 21534 25284 21586
rect 25228 21028 25284 21534
rect 25340 21588 25396 21598
rect 25340 21494 25396 21532
rect 25452 21586 25508 21598
rect 25452 21534 25454 21586
rect 25506 21534 25508 21586
rect 25228 20962 25284 20972
rect 25340 20804 25396 20814
rect 25340 20710 25396 20748
rect 25452 20580 25508 21534
rect 25228 20524 25508 20580
rect 25228 20020 25284 20524
rect 25228 19954 25284 19964
rect 25340 20244 25396 20254
rect 25340 20018 25396 20188
rect 25564 20130 25620 23436
rect 25676 23156 25732 23166
rect 25676 23062 25732 23100
rect 25788 21586 25844 23884
rect 25900 22596 25956 23996
rect 26348 23938 26404 23950
rect 26348 23886 26350 23938
rect 26402 23886 26404 23938
rect 26124 23826 26180 23838
rect 26124 23774 26126 23826
rect 26178 23774 26180 23826
rect 26012 23268 26068 23278
rect 26124 23268 26180 23774
rect 26012 23266 26180 23268
rect 26012 23214 26014 23266
rect 26066 23214 26180 23266
rect 26012 23212 26180 23214
rect 26348 23266 26404 23886
rect 26460 23380 26516 24446
rect 26460 23314 26516 23324
rect 26348 23214 26350 23266
rect 26402 23214 26404 23266
rect 26012 23202 26068 23212
rect 26348 23202 26404 23214
rect 26572 22820 26628 24556
rect 26908 24612 26964 24622
rect 26908 24518 26964 24556
rect 27132 23714 27188 23726
rect 27132 23662 27134 23714
rect 27186 23662 27188 23714
rect 26684 23268 26740 23278
rect 26684 23156 26740 23212
rect 26684 23154 26852 23156
rect 26684 23102 26686 23154
rect 26738 23102 26852 23154
rect 26684 23100 26852 23102
rect 26684 23090 26740 23100
rect 26572 22754 26628 22764
rect 26572 22596 26628 22606
rect 25900 22540 26068 22596
rect 25900 22370 25956 22382
rect 25900 22318 25902 22370
rect 25954 22318 25956 22370
rect 25900 21924 25956 22318
rect 26012 22036 26068 22540
rect 26572 22502 26628 22540
rect 26124 22372 26180 22382
rect 26460 22372 26516 22410
rect 26124 22370 26292 22372
rect 26124 22318 26126 22370
rect 26178 22318 26292 22370
rect 26124 22316 26292 22318
rect 26124 22306 26180 22316
rect 26236 22260 26292 22316
rect 26460 22306 26516 22316
rect 26684 22372 26740 22382
rect 26684 22278 26740 22316
rect 26236 22204 26404 22260
rect 26348 22148 26404 22204
rect 26796 22148 26852 23100
rect 26908 23042 26964 23054
rect 26908 22990 26910 23042
rect 26962 22990 26964 23042
rect 26908 22708 26964 22990
rect 26908 22642 26964 22652
rect 27020 22372 27076 22382
rect 27020 22278 27076 22316
rect 26348 22092 26852 22148
rect 26012 21980 26404 22036
rect 25900 21858 25956 21868
rect 26012 21812 26068 21822
rect 26012 21718 26068 21756
rect 26236 21700 26292 21738
rect 26236 21634 26292 21644
rect 25788 21534 25790 21586
rect 25842 21534 25844 21586
rect 25564 20078 25566 20130
rect 25618 20078 25620 20130
rect 25564 20066 25620 20078
rect 25676 20916 25732 20926
rect 25340 19966 25342 20018
rect 25394 19966 25396 20018
rect 25340 19954 25396 19966
rect 25452 19796 25508 19806
rect 25116 19348 25172 19358
rect 25116 19254 25172 19292
rect 24556 18274 24612 18284
rect 24668 19180 25060 19236
rect 24668 18674 24724 19180
rect 24668 18622 24670 18674
rect 24722 18622 24724 18674
rect 24556 17108 24612 17118
rect 24444 17052 24556 17108
rect 24332 16882 24388 17052
rect 24332 16830 24334 16882
rect 24386 16830 24388 16882
rect 24332 16818 24388 16830
rect 23884 16034 23940 16044
rect 23996 16098 24052 16110
rect 23996 16046 23998 16098
rect 24050 16046 24052 16098
rect 23884 15874 23940 15886
rect 23884 15822 23886 15874
rect 23938 15822 23940 15874
rect 23772 15316 23828 15326
rect 23884 15316 23940 15822
rect 23996 15876 24052 16046
rect 24444 15876 24500 15886
rect 23996 15810 24052 15820
rect 24220 15820 24444 15876
rect 23772 15314 23940 15316
rect 23772 15262 23774 15314
rect 23826 15262 23940 15314
rect 23772 15260 23940 15262
rect 23772 15250 23828 15260
rect 24220 15202 24276 15820
rect 24444 15810 24500 15820
rect 24220 15150 24222 15202
rect 24274 15150 24276 15202
rect 24220 15148 24276 15150
rect 24444 15540 24500 15550
rect 23548 15092 23604 15102
rect 24220 15092 24388 15148
rect 23548 14530 23604 15036
rect 24108 14756 24164 14766
rect 23548 14478 23550 14530
rect 23602 14478 23604 14530
rect 23548 14466 23604 14478
rect 23996 14532 24052 14542
rect 24108 14532 24164 14700
rect 23996 14530 24164 14532
rect 23996 14478 23998 14530
rect 24050 14478 24164 14530
rect 23996 14476 24164 14478
rect 24332 14530 24388 15092
rect 24332 14478 24334 14530
rect 24386 14478 24388 14530
rect 23996 14466 24052 14476
rect 22988 14420 23044 14430
rect 22876 14418 23044 14420
rect 22876 14366 22990 14418
rect 23042 14366 23044 14418
rect 22876 14364 23044 14366
rect 22988 14196 23044 14364
rect 23100 14420 23156 14430
rect 23100 14308 23156 14364
rect 23660 14420 23716 14430
rect 23324 14308 23380 14318
rect 23100 14306 23380 14308
rect 23100 14254 23326 14306
rect 23378 14254 23380 14306
rect 23100 14252 23380 14254
rect 23324 14242 23380 14252
rect 23436 14308 23492 14318
rect 23660 14308 23716 14364
rect 23436 14306 23716 14308
rect 23436 14254 23438 14306
rect 23490 14254 23716 14306
rect 23436 14252 23716 14254
rect 23436 14242 23492 14252
rect 22988 14140 23156 14196
rect 23100 13858 23156 14140
rect 23100 13806 23102 13858
rect 23154 13806 23156 13858
rect 23100 13794 23156 13806
rect 23324 13972 23380 13982
rect 22988 13748 23044 13758
rect 22988 13654 23044 13692
rect 22764 13634 22820 13646
rect 22764 13582 22766 13634
rect 22818 13582 22820 13634
rect 22764 13524 22820 13582
rect 22764 13458 22820 13468
rect 22540 12402 22708 12404
rect 22540 12350 22542 12402
rect 22594 12350 22708 12402
rect 22540 12348 22708 12350
rect 22764 13300 22820 13310
rect 22764 12402 22820 13244
rect 22764 12350 22766 12402
rect 22818 12350 22820 12402
rect 22540 12338 22596 12348
rect 22764 12292 22820 12350
rect 23100 13300 23156 13310
rect 23100 12402 23156 13244
rect 23100 12350 23102 12402
rect 23154 12350 23156 12402
rect 23100 12338 23156 12350
rect 22764 12236 23044 12292
rect 22428 12180 22484 12190
rect 22428 9492 22484 12124
rect 22652 12180 22708 12190
rect 22652 11956 22708 12124
rect 22652 11890 22708 11900
rect 22876 11956 22932 11966
rect 22540 11620 22596 11630
rect 22540 11394 22596 11564
rect 22764 11620 22820 11630
rect 22876 11620 22932 11900
rect 22764 11618 22932 11620
rect 22764 11566 22766 11618
rect 22818 11566 22932 11618
rect 22764 11564 22932 11566
rect 22988 11620 23044 12236
rect 22764 11554 22820 11564
rect 22988 11554 23044 11564
rect 23212 12180 23268 12190
rect 22988 11396 23044 11406
rect 22540 11342 22542 11394
rect 22594 11342 22596 11394
rect 22540 11330 22596 11342
rect 22876 11394 23044 11396
rect 22876 11342 22990 11394
rect 23042 11342 23044 11394
rect 22876 11340 23044 11342
rect 22540 10724 22596 10734
rect 22540 10630 22596 10668
rect 22764 10388 22820 10398
rect 22764 9826 22820 10332
rect 22764 9774 22766 9826
rect 22818 9774 22820 9826
rect 22764 9762 22820 9774
rect 22540 9716 22596 9726
rect 22540 9622 22596 9660
rect 22652 9604 22708 9614
rect 22652 9510 22708 9548
rect 22428 9426 22484 9436
rect 22764 9492 22820 9502
rect 22764 9042 22820 9436
rect 22764 8990 22766 9042
rect 22818 8990 22820 9042
rect 22764 8978 22820 8990
rect 22316 8418 22372 8428
rect 22428 8596 22484 8606
rect 22428 7250 22484 8540
rect 22876 7924 22932 11340
rect 22988 11330 23044 11340
rect 23100 11396 23156 11406
rect 23100 11302 23156 11340
rect 22988 10836 23044 10846
rect 22988 10742 23044 10780
rect 23212 10612 23268 12124
rect 22876 7858 22932 7868
rect 22988 10556 23268 10612
rect 22540 7700 22596 7710
rect 22988 7700 23044 10556
rect 23100 10388 23156 10398
rect 23324 10388 23380 13916
rect 23548 13972 23604 13982
rect 23604 13916 23716 13972
rect 23548 13906 23604 13916
rect 23548 13524 23604 13534
rect 23548 12962 23604 13468
rect 23548 12910 23550 12962
rect 23602 12910 23604 12962
rect 23548 12898 23604 12910
rect 23436 11620 23492 11630
rect 23436 10836 23492 11564
rect 23548 11620 23604 11630
rect 23660 11620 23716 13916
rect 23772 13860 23828 13870
rect 23772 13746 23828 13804
rect 23772 13694 23774 13746
rect 23826 13694 23828 13746
rect 23772 13682 23828 13694
rect 23996 13860 24052 13870
rect 24332 13860 24388 14478
rect 23996 13858 24388 13860
rect 23996 13806 23998 13858
rect 24050 13806 24388 13858
rect 23996 13804 24388 13806
rect 24444 13858 24500 15484
rect 24444 13806 24446 13858
rect 24498 13806 24500 13858
rect 23884 13300 23940 13310
rect 23996 13300 24052 13804
rect 24444 13748 24500 13806
rect 23940 13244 24052 13300
rect 24108 13692 24500 13748
rect 23884 13234 23940 13244
rect 23772 12066 23828 12078
rect 23772 12014 23774 12066
rect 23826 12014 23828 12066
rect 23772 11844 23828 12014
rect 23772 11778 23828 11788
rect 23548 11618 23716 11620
rect 23548 11566 23550 11618
rect 23602 11566 23716 11618
rect 23548 11564 23716 11566
rect 23548 11554 23604 11564
rect 23772 11396 23828 11406
rect 23772 11302 23828 11340
rect 23996 11394 24052 11406
rect 23996 11342 23998 11394
rect 24050 11342 24052 11394
rect 23884 11172 23940 11182
rect 23548 10836 23604 10846
rect 23436 10834 23604 10836
rect 23436 10782 23550 10834
rect 23602 10782 23604 10834
rect 23436 10780 23604 10782
rect 23324 10332 23492 10388
rect 23100 9268 23156 10332
rect 23436 10164 23492 10332
rect 23324 10052 23380 10062
rect 23324 9938 23380 9996
rect 23324 9886 23326 9938
rect 23378 9886 23380 9938
rect 23324 9874 23380 9886
rect 23436 9826 23492 10108
rect 23436 9774 23438 9826
rect 23490 9774 23492 9826
rect 23436 9762 23492 9774
rect 23212 9602 23268 9614
rect 23548 9604 23604 10780
rect 23772 10724 23828 10734
rect 23772 10610 23828 10668
rect 23772 10558 23774 10610
rect 23826 10558 23828 10610
rect 23772 10546 23828 10558
rect 23212 9550 23214 9602
rect 23266 9550 23268 9602
rect 23212 9492 23268 9550
rect 23436 9548 23604 9604
rect 23772 9826 23828 9838
rect 23772 9774 23774 9826
rect 23826 9774 23828 9826
rect 23212 9436 23380 9492
rect 23212 9268 23268 9278
rect 23100 9266 23268 9268
rect 23100 9214 23214 9266
rect 23266 9214 23268 9266
rect 23100 9212 23268 9214
rect 23212 9202 23268 9212
rect 23324 8932 23380 9436
rect 22540 7698 23044 7700
rect 22540 7646 22542 7698
rect 22594 7646 22990 7698
rect 23042 7646 23044 7698
rect 22540 7644 23044 7646
rect 22540 7634 22596 7644
rect 22988 7634 23044 7644
rect 23100 8820 23156 8830
rect 23100 7476 23156 8764
rect 23324 8708 23380 8876
rect 22428 7198 22430 7250
rect 22482 7198 22484 7250
rect 22428 7186 22484 7198
rect 22652 7420 23156 7476
rect 23212 8652 23380 8708
rect 22204 6962 22260 6972
rect 21980 6860 22148 6916
rect 21980 6468 22036 6860
rect 22092 6692 22148 6702
rect 22652 6692 22708 7420
rect 22148 6636 22260 6692
rect 22092 6626 22148 6636
rect 22092 6468 22148 6478
rect 21980 6466 22148 6468
rect 21980 6414 22094 6466
rect 22146 6414 22148 6466
rect 21980 6412 22148 6414
rect 22092 6402 22148 6412
rect 22092 6132 22148 6142
rect 22204 6132 22260 6636
rect 22540 6690 22708 6692
rect 22540 6638 22654 6690
rect 22706 6638 22708 6690
rect 22540 6636 22708 6638
rect 22092 6130 22260 6132
rect 22092 6078 22094 6130
rect 22146 6078 22260 6130
rect 22092 6076 22260 6078
rect 22316 6466 22372 6478
rect 22316 6414 22318 6466
rect 22370 6414 22372 6466
rect 22092 6066 22148 6076
rect 22316 5908 22372 6414
rect 21756 5070 21758 5122
rect 21810 5070 21812 5122
rect 21756 5058 21812 5070
rect 21980 5122 22036 5134
rect 21980 5070 21982 5122
rect 22034 5070 22036 5122
rect 21084 4562 21364 4564
rect 21084 4510 21086 4562
rect 21138 4510 21364 4562
rect 21084 4508 21364 4510
rect 21420 5010 21476 5022
rect 21420 4958 21422 5010
rect 21474 4958 21476 5010
rect 21420 4564 21476 4958
rect 21084 4498 21140 4508
rect 21420 4498 21476 4508
rect 21532 4898 21588 4910
rect 21532 4846 21534 4898
rect 21586 4846 21588 4898
rect 21532 4452 21588 4846
rect 21980 4676 22036 5070
rect 22204 5124 22260 5134
rect 22204 5030 22260 5068
rect 22316 5012 22372 5852
rect 22428 6468 22484 6478
rect 22428 5234 22484 6412
rect 22428 5182 22430 5234
rect 22482 5182 22484 5234
rect 22428 5170 22484 5182
rect 22316 4956 22484 5012
rect 21980 4620 22372 4676
rect 21868 4564 21924 4574
rect 21868 4470 21924 4508
rect 21532 4386 21588 4396
rect 22204 4452 22260 4462
rect 22204 4358 22260 4396
rect 21532 4226 21588 4238
rect 21532 4174 21534 4226
rect 21586 4174 21588 4226
rect 21532 4004 21588 4174
rect 22316 4114 22372 4620
rect 22428 4450 22484 4956
rect 22428 4398 22430 4450
rect 22482 4398 22484 4450
rect 22428 4386 22484 4398
rect 22316 4062 22318 4114
rect 22370 4062 22372 4114
rect 22316 4050 22372 4062
rect 21532 3938 21588 3948
rect 22540 3892 22596 6636
rect 22652 6626 22708 6636
rect 23100 7250 23156 7262
rect 23100 7198 23102 7250
rect 23154 7198 23156 7250
rect 23100 6802 23156 7198
rect 23100 6750 23102 6802
rect 23154 6750 23156 6802
rect 22652 6020 22708 6030
rect 22652 5926 22708 5964
rect 22988 5908 23044 5918
rect 22988 5814 23044 5852
rect 22764 5794 22820 5806
rect 22764 5742 22766 5794
rect 22818 5742 22820 5794
rect 22652 5124 22708 5134
rect 22764 5124 22820 5742
rect 23100 5684 23156 6750
rect 23100 5618 23156 5628
rect 22652 5122 22820 5124
rect 22652 5070 22654 5122
rect 22706 5070 22820 5122
rect 22652 5068 22820 5070
rect 23212 5124 23268 8652
rect 23324 8484 23380 8494
rect 23324 8258 23380 8428
rect 23324 8206 23326 8258
rect 23378 8206 23380 8258
rect 23324 8194 23380 8206
rect 23436 7924 23492 9548
rect 23772 9492 23828 9774
rect 22652 5058 22708 5068
rect 23212 5058 23268 5068
rect 23324 7868 23492 7924
rect 23548 9436 23772 9492
rect 23324 6130 23380 7868
rect 23436 7700 23492 7710
rect 23548 7700 23604 9436
rect 23772 9398 23828 9436
rect 23884 9156 23940 11116
rect 23884 9090 23940 9100
rect 23996 8484 24052 11342
rect 24108 11396 24164 13692
rect 24220 13076 24276 13086
rect 24220 12402 24276 13020
rect 24220 12350 24222 12402
rect 24274 12350 24276 12402
rect 24220 12338 24276 12350
rect 24444 12516 24500 12526
rect 24444 12290 24500 12460
rect 24444 12238 24446 12290
rect 24498 12238 24500 12290
rect 24444 12226 24500 12238
rect 24332 12066 24388 12078
rect 24332 12014 24334 12066
rect 24386 12014 24388 12066
rect 24108 11330 24164 11340
rect 24220 11956 24276 11966
rect 24332 11956 24388 12014
rect 24556 11956 24612 17052
rect 24668 16996 24724 18622
rect 25004 19010 25060 19022
rect 25004 18958 25006 19010
rect 25058 18958 25060 19010
rect 25004 18676 25060 18958
rect 25004 18610 25060 18620
rect 25228 19012 25284 19022
rect 25228 18452 25284 18956
rect 25452 19012 25508 19740
rect 25676 19572 25732 20860
rect 25788 19796 25844 21534
rect 26348 21586 26404 21980
rect 26348 21534 26350 21586
rect 26402 21534 26404 21586
rect 26236 21140 26292 21150
rect 26236 20804 26292 21084
rect 26124 20802 26292 20804
rect 26124 20750 26238 20802
rect 26290 20750 26292 20802
rect 26124 20748 26292 20750
rect 26012 20692 26068 20702
rect 26012 20598 26068 20636
rect 26012 19908 26068 19918
rect 26012 19814 26068 19852
rect 25788 19730 25844 19740
rect 25676 19506 25732 19516
rect 25452 18946 25508 18956
rect 25676 19234 25732 19246
rect 25676 19182 25678 19234
rect 25730 19182 25732 19234
rect 25676 19124 25732 19182
rect 26012 19236 26068 19246
rect 26012 19142 26068 19180
rect 25900 19124 25956 19134
rect 25676 19122 25956 19124
rect 25676 19070 25902 19122
rect 25954 19070 25956 19122
rect 25676 19068 25956 19070
rect 25452 18452 25508 18462
rect 25228 18450 25508 18452
rect 25228 18398 25454 18450
rect 25506 18398 25508 18450
rect 25228 18396 25508 18398
rect 25452 18386 25508 18396
rect 25564 18338 25620 18350
rect 25564 18286 25566 18338
rect 25618 18286 25620 18338
rect 25564 18228 25620 18286
rect 25004 18116 25060 18126
rect 25060 18060 25172 18116
rect 25004 18050 25060 18060
rect 24780 17778 24836 17790
rect 24780 17726 24782 17778
rect 24834 17726 24836 17778
rect 24780 17106 24836 17726
rect 24780 17054 24782 17106
rect 24834 17054 24836 17106
rect 24780 17042 24836 17054
rect 24668 16930 24724 16940
rect 25116 16772 25172 18060
rect 25452 17780 25508 17790
rect 25452 17108 25508 17724
rect 25340 17106 25508 17108
rect 25340 17054 25454 17106
rect 25506 17054 25508 17106
rect 25340 17052 25508 17054
rect 25228 16772 25284 16782
rect 25116 16770 25284 16772
rect 25116 16718 25230 16770
rect 25282 16718 25284 16770
rect 25116 16716 25284 16718
rect 25228 16706 25284 16716
rect 25340 16324 25396 17052
rect 25452 17042 25508 17052
rect 25340 16258 25396 16268
rect 25452 16770 25508 16782
rect 25452 16718 25454 16770
rect 25506 16718 25508 16770
rect 25004 16156 25284 16212
rect 25004 16100 25060 16156
rect 25004 16006 25060 16044
rect 25116 15986 25172 15998
rect 25116 15934 25118 15986
rect 25170 15934 25172 15986
rect 25116 15876 25172 15934
rect 25116 15810 25172 15820
rect 24668 15428 24724 15438
rect 24668 15334 24724 15372
rect 24892 15204 24948 15214
rect 24780 14418 24836 14430
rect 24780 14366 24782 14418
rect 24834 14366 24836 14418
rect 24780 13860 24836 14366
rect 24780 13794 24836 13804
rect 24892 12962 24948 15148
rect 25228 15148 25284 16156
rect 25228 15092 25396 15148
rect 25116 14868 25172 14878
rect 25172 14812 25284 14868
rect 25004 14530 25060 14542
rect 25004 14478 25006 14530
rect 25058 14478 25060 14530
rect 25004 14308 25060 14478
rect 25004 14242 25060 14252
rect 25116 13412 25172 14812
rect 25228 14530 25284 14812
rect 25228 14478 25230 14530
rect 25282 14478 25284 14530
rect 25228 14466 25284 14478
rect 25228 13972 25284 13982
rect 25340 13972 25396 15092
rect 25228 13970 25396 13972
rect 25228 13918 25230 13970
rect 25282 13918 25396 13970
rect 25228 13916 25396 13918
rect 25228 13906 25284 13916
rect 25452 13748 25508 16718
rect 25564 16212 25620 18172
rect 25564 16146 25620 16156
rect 25676 15988 25732 19068
rect 25900 19058 25956 19068
rect 25900 18340 25956 18350
rect 25900 17780 25956 18284
rect 25900 17666 25956 17724
rect 25900 17614 25902 17666
rect 25954 17614 25956 17666
rect 25900 17602 25956 17614
rect 26012 18338 26068 18350
rect 26012 18286 26014 18338
rect 26066 18286 26068 18338
rect 26012 17668 26068 18286
rect 26012 17602 26068 17612
rect 25788 16996 25844 17006
rect 25788 16882 25844 16940
rect 25788 16830 25790 16882
rect 25842 16830 25844 16882
rect 25788 16818 25844 16830
rect 25900 16098 25956 16110
rect 25900 16046 25902 16098
rect 25954 16046 25956 16098
rect 25564 15932 25732 15988
rect 25788 15986 25844 15998
rect 25788 15934 25790 15986
rect 25842 15934 25844 15986
rect 25564 14756 25620 15932
rect 25788 15652 25844 15934
rect 25788 15586 25844 15596
rect 25788 15314 25844 15326
rect 25788 15262 25790 15314
rect 25842 15262 25844 15314
rect 25676 15204 25732 15242
rect 25676 15138 25732 15148
rect 25676 14756 25732 14766
rect 25564 14700 25676 14756
rect 24892 12910 24894 12962
rect 24946 12910 24948 12962
rect 24892 12898 24948 12910
rect 25004 13356 25172 13412
rect 25340 13692 25508 13748
rect 25564 13858 25620 13870
rect 25564 13806 25566 13858
rect 25618 13806 25620 13858
rect 24332 11900 24500 11956
rect 24220 11394 24276 11900
rect 24332 11732 24388 11742
rect 24332 11506 24388 11676
rect 24332 11454 24334 11506
rect 24386 11454 24388 11506
rect 24332 11442 24388 11454
rect 24220 11342 24222 11394
rect 24274 11342 24276 11394
rect 24220 11330 24276 11342
rect 24444 11282 24500 11900
rect 24556 11890 24612 11900
rect 24892 11732 24948 11742
rect 24892 11618 24948 11676
rect 24892 11566 24894 11618
rect 24946 11566 24948 11618
rect 24892 11554 24948 11566
rect 25004 11620 25060 13356
rect 25116 13188 25172 13198
rect 25116 13094 25172 13132
rect 25228 13074 25284 13086
rect 25228 13022 25230 13074
rect 25282 13022 25284 13074
rect 25004 11554 25060 11564
rect 25116 11844 25172 11854
rect 24444 11230 24446 11282
rect 24498 11230 24500 11282
rect 24332 11172 24388 11182
rect 24444 11172 24500 11230
rect 25004 11394 25060 11406
rect 25004 11342 25006 11394
rect 25058 11342 25060 11394
rect 24388 11116 24500 11172
rect 24556 11172 24612 11182
rect 24332 11106 24388 11116
rect 24108 10836 24164 10846
rect 24108 10742 24164 10780
rect 24332 10836 24388 10846
rect 24332 10742 24388 10780
rect 24444 10836 24500 10846
rect 24556 10836 24612 11116
rect 24444 10834 24612 10836
rect 24444 10782 24446 10834
rect 24498 10782 24612 10834
rect 24444 10780 24612 10782
rect 25004 10836 25060 11342
rect 24444 10770 24500 10780
rect 25004 10770 25060 10780
rect 24444 10164 24500 10174
rect 24108 10052 24164 10062
rect 24108 9826 24164 9996
rect 24108 9774 24110 9826
rect 24162 9774 24164 9826
rect 24108 9762 24164 9774
rect 24220 9828 24276 9838
rect 24220 9714 24276 9772
rect 24444 9826 24500 10108
rect 24444 9774 24446 9826
rect 24498 9774 24500 9826
rect 24444 9762 24500 9774
rect 24220 9662 24222 9714
rect 24274 9662 24276 9714
rect 24220 9650 24276 9662
rect 25116 9602 25172 11788
rect 25116 9550 25118 9602
rect 25170 9550 25172 9602
rect 24108 9380 24164 9390
rect 24108 9268 24164 9324
rect 24108 9266 24276 9268
rect 24108 9214 24110 9266
rect 24162 9214 24276 9266
rect 24108 9212 24276 9214
rect 24108 9202 24164 9212
rect 23996 8428 24164 8484
rect 23772 8258 23828 8270
rect 23772 8206 23774 8258
rect 23826 8206 23828 8258
rect 23772 8148 23828 8206
rect 23772 8082 23828 8092
rect 23996 8258 24052 8270
rect 23996 8206 23998 8258
rect 24050 8206 24052 8258
rect 23436 7698 23604 7700
rect 23436 7646 23438 7698
rect 23490 7646 23604 7698
rect 23436 7644 23604 7646
rect 23660 7924 23716 7934
rect 23436 7634 23492 7644
rect 23324 6078 23326 6130
rect 23378 6078 23380 6130
rect 22764 4900 22820 4910
rect 22764 4806 22820 4844
rect 22876 4898 22932 4910
rect 22876 4846 22878 4898
rect 22930 4846 22932 4898
rect 22876 4788 22932 4846
rect 22764 4676 22820 4686
rect 22764 4338 22820 4620
rect 22876 4452 22932 4732
rect 23324 4564 23380 6078
rect 23660 6356 23716 7868
rect 23884 7700 23940 7710
rect 23884 7606 23940 7644
rect 23996 7364 24052 8206
rect 24108 7476 24164 8428
rect 24108 7410 24164 7420
rect 24220 7474 24276 9212
rect 24556 9156 24612 9166
rect 24556 9062 24612 9100
rect 24444 9044 24500 9054
rect 24444 8950 24500 8988
rect 24780 9044 24836 9054
rect 24780 8950 24836 8988
rect 25004 8484 25060 8494
rect 25004 8390 25060 8428
rect 24892 8372 24948 8382
rect 24892 8258 24948 8316
rect 24892 8206 24894 8258
rect 24946 8206 24948 8258
rect 24220 7422 24222 7474
rect 24274 7422 24276 7474
rect 23996 7298 24052 7308
rect 24220 7364 24276 7422
rect 24556 7924 24612 7934
rect 24556 7474 24612 7868
rect 24556 7422 24558 7474
rect 24610 7422 24612 7474
rect 24556 7410 24612 7422
rect 24220 7298 24276 7308
rect 24668 7364 24724 7374
rect 24668 7270 24724 7308
rect 23884 7252 23940 7262
rect 23660 6130 23716 6300
rect 23660 6078 23662 6130
rect 23714 6078 23716 6130
rect 23660 6066 23716 6078
rect 23772 6468 23828 6478
rect 23324 4452 23380 4508
rect 23772 5908 23828 6412
rect 23772 4564 23828 5852
rect 23884 5234 23940 7196
rect 24332 7252 24388 7262
rect 24556 7252 24612 7262
rect 24332 7250 24500 7252
rect 24332 7198 24334 7250
rect 24386 7198 24500 7250
rect 24332 7196 24500 7198
rect 24332 7186 24388 7196
rect 24108 6804 24164 6814
rect 23996 6748 24108 6804
rect 23996 6690 24052 6748
rect 24108 6738 24164 6748
rect 24444 6804 24500 7196
rect 24444 6738 24500 6748
rect 23996 6638 23998 6690
rect 24050 6638 24052 6690
rect 23996 6626 24052 6638
rect 24108 6580 24164 6590
rect 24108 5460 24164 6524
rect 24444 6580 24500 6590
rect 24556 6580 24612 7196
rect 24892 7252 24948 8206
rect 24892 7186 24948 7196
rect 25004 8148 25060 8158
rect 24892 7028 24948 7038
rect 24892 6802 24948 6972
rect 25004 6914 25060 8092
rect 25004 6862 25006 6914
rect 25058 6862 25060 6914
rect 25004 6850 25060 6862
rect 24892 6750 24894 6802
rect 24946 6750 24948 6802
rect 24892 6738 24948 6750
rect 24500 6524 24612 6580
rect 24668 6690 24724 6702
rect 24668 6638 24670 6690
rect 24722 6638 24724 6690
rect 24444 6486 24500 6524
rect 24668 6468 24724 6638
rect 24668 6402 24724 6412
rect 24332 6020 24388 6030
rect 24332 5926 24388 5964
rect 24780 6020 24836 6030
rect 24780 5926 24836 5964
rect 25116 5684 25172 9550
rect 25228 10386 25284 13022
rect 25340 10724 25396 13692
rect 25452 13524 25508 13534
rect 25452 12402 25508 13468
rect 25452 12350 25454 12402
rect 25506 12350 25508 12402
rect 25452 12338 25508 12350
rect 25564 12516 25620 13806
rect 25676 13076 25732 14700
rect 25676 13010 25732 13020
rect 25452 11620 25508 11630
rect 25452 11284 25508 11564
rect 25452 11218 25508 11228
rect 25340 10658 25396 10668
rect 25228 10334 25230 10386
rect 25282 10334 25284 10386
rect 25228 8372 25284 10334
rect 25340 10498 25396 10510
rect 25340 10446 25342 10498
rect 25394 10446 25396 10498
rect 25340 9716 25396 10446
rect 25452 10052 25508 10062
rect 25452 9958 25508 9996
rect 25340 8708 25396 9660
rect 25564 9604 25620 12460
rect 25788 11844 25844 15262
rect 25900 15092 25956 16046
rect 25900 13970 25956 15036
rect 26124 14420 26180 20748
rect 26236 20738 26292 20748
rect 26348 20356 26404 21534
rect 26796 21810 26852 22092
rect 26908 21924 26964 21934
rect 27132 21924 27188 23662
rect 27356 22148 27412 26012
rect 27468 25396 27524 27804
rect 27580 27186 27636 28028
rect 27692 27990 27748 28028
rect 27804 27748 27860 30268
rect 27916 29988 27972 29998
rect 27916 29894 27972 29932
rect 28140 29426 28196 31276
rect 30044 31332 30100 31726
rect 30044 31266 30100 31276
rect 28140 29374 28142 29426
rect 28194 29374 28196 29426
rect 28140 29362 28196 29374
rect 28476 29986 28532 29998
rect 28476 29934 28478 29986
rect 28530 29934 28532 29986
rect 28476 28644 28532 29934
rect 30268 29876 30324 29886
rect 30380 29876 30436 33964
rect 31052 33954 31108 33966
rect 30828 32564 30884 32574
rect 30884 32508 30996 32564
rect 30828 32498 30884 32508
rect 30604 32452 30660 32462
rect 30604 31892 30660 32396
rect 30828 32004 30884 32014
rect 30828 31892 30884 31948
rect 30604 31836 30884 31892
rect 30492 31780 30548 31790
rect 30492 31778 30772 31780
rect 30492 31726 30494 31778
rect 30546 31726 30772 31778
rect 30492 31724 30772 31726
rect 30492 31714 30548 31724
rect 30716 30098 30772 31724
rect 30716 30046 30718 30098
rect 30770 30046 30772 30098
rect 30716 30034 30772 30046
rect 30324 29820 30436 29876
rect 30828 29988 30884 31836
rect 30268 29810 30324 29820
rect 30828 29650 30884 29932
rect 30828 29598 30830 29650
rect 30882 29598 30884 29650
rect 30828 29586 30884 29598
rect 28588 29428 28644 29438
rect 28588 29334 28644 29372
rect 29148 29428 29204 29438
rect 28476 28588 28644 28644
rect 28476 28418 28532 28430
rect 28476 28366 28478 28418
rect 28530 28366 28532 28418
rect 28476 27972 28532 28366
rect 28588 28084 28644 28588
rect 29148 28530 29204 29372
rect 29484 28644 29540 28654
rect 29484 28550 29540 28588
rect 29148 28478 29150 28530
rect 29202 28478 29204 28530
rect 29148 28466 29204 28478
rect 28588 28018 28644 28028
rect 29036 28084 29092 28094
rect 29820 28084 29876 28094
rect 30828 28084 30884 28094
rect 30940 28084 30996 32508
rect 31836 31332 31892 31342
rect 31836 31106 31892 31276
rect 31836 31054 31838 31106
rect 31890 31054 31892 31106
rect 31836 31042 31892 31054
rect 31948 31108 32004 31118
rect 31836 30212 31892 30222
rect 31052 30100 31108 30110
rect 31724 30100 31780 30110
rect 31052 30098 31780 30100
rect 31052 30046 31054 30098
rect 31106 30046 31726 30098
rect 31778 30046 31780 30098
rect 31052 30044 31780 30046
rect 31052 30034 31108 30044
rect 31724 30034 31780 30044
rect 31836 29876 31892 30156
rect 31948 29988 32004 31052
rect 32060 30322 32116 30334
rect 32060 30270 32062 30322
rect 32114 30270 32116 30322
rect 32060 30212 32116 30270
rect 32060 30146 32116 30156
rect 31948 29932 32116 29988
rect 31388 29820 31892 29876
rect 31388 28866 31444 29820
rect 31612 29652 31668 29662
rect 31612 29558 31668 29596
rect 31724 29650 31780 29662
rect 31724 29598 31726 29650
rect 31778 29598 31780 29650
rect 31388 28814 31390 28866
rect 31442 28814 31444 28866
rect 31388 28802 31444 28814
rect 31052 28644 31108 28654
rect 31724 28644 31780 29598
rect 31948 29538 32004 29550
rect 31948 29486 31950 29538
rect 32002 29486 32004 29538
rect 31948 29316 32004 29486
rect 32060 29538 32116 29932
rect 32060 29486 32062 29538
rect 32114 29486 32116 29538
rect 32060 29474 32116 29486
rect 32172 29652 32228 29662
rect 31948 29260 32116 29316
rect 31948 28756 32004 28766
rect 32060 28756 32116 29260
rect 32004 28700 32116 28756
rect 31948 28690 32004 28700
rect 31836 28644 31892 28654
rect 31724 28642 31892 28644
rect 31724 28590 31838 28642
rect 31890 28590 31892 28642
rect 31724 28588 31892 28590
rect 31052 28550 31108 28588
rect 31836 28578 31892 28588
rect 32172 28530 32228 29596
rect 32172 28478 32174 28530
rect 32226 28478 32228 28530
rect 32172 28466 32228 28478
rect 29092 28028 29316 28084
rect 29036 27990 29092 28028
rect 28140 27916 28532 27972
rect 27804 27682 27860 27692
rect 28028 27858 28084 27870
rect 28028 27806 28030 27858
rect 28082 27806 28084 27858
rect 27692 27300 27748 27310
rect 28028 27300 28084 27806
rect 27692 27298 28084 27300
rect 27692 27246 27694 27298
rect 27746 27246 28084 27298
rect 27692 27244 28084 27246
rect 27692 27234 27748 27244
rect 27580 27134 27582 27186
rect 27634 27134 27636 27186
rect 27580 27122 27636 27134
rect 27804 27076 27860 27086
rect 27692 26402 27748 26414
rect 27692 26350 27694 26402
rect 27746 26350 27748 26402
rect 27580 25396 27636 25406
rect 27468 25340 27580 25396
rect 27580 25330 27636 25340
rect 27692 25284 27748 26350
rect 27468 24948 27524 24958
rect 27692 24948 27748 25228
rect 27468 24946 27748 24948
rect 27468 24894 27470 24946
rect 27522 24894 27748 24946
rect 27468 24892 27748 24894
rect 27804 24946 27860 27020
rect 28028 27074 28084 27244
rect 28028 27022 28030 27074
rect 28082 27022 28084 27074
rect 28028 27010 28084 27022
rect 28140 26852 28196 27916
rect 27916 26796 28196 26852
rect 28252 27748 28308 27758
rect 27916 25956 27972 26796
rect 28252 26628 28308 27692
rect 28476 27746 28532 27758
rect 28476 27694 28478 27746
rect 28530 27694 28532 27746
rect 28476 27524 28532 27694
rect 28476 27458 28532 27468
rect 28924 27636 28980 27646
rect 28476 27186 28532 27198
rect 28476 27134 28478 27186
rect 28530 27134 28532 27186
rect 28476 26908 28532 27134
rect 28476 26852 28644 26908
rect 27916 25890 27972 25900
rect 28028 26572 28308 26628
rect 27804 24894 27806 24946
rect 27858 24894 27860 24946
rect 27468 24882 27524 24892
rect 27468 23940 27524 23950
rect 27804 23940 27860 24894
rect 27468 23938 27860 23940
rect 27468 23886 27470 23938
rect 27522 23886 27860 23938
rect 27468 23884 27860 23886
rect 27916 25396 27972 25406
rect 27468 23874 27524 23884
rect 27468 23268 27524 23278
rect 27468 23154 27524 23212
rect 27468 23102 27470 23154
rect 27522 23102 27524 23154
rect 27468 23090 27524 23102
rect 27580 23156 27636 23166
rect 27580 22370 27636 23100
rect 27580 22318 27582 22370
rect 27634 22318 27636 22370
rect 27580 22306 27636 22318
rect 27356 22092 27860 22148
rect 26964 21868 27076 21924
rect 27132 21868 27524 21924
rect 26908 21858 26964 21868
rect 26796 21758 26798 21810
rect 26850 21758 26852 21810
rect 26796 21476 26852 21758
rect 26796 21410 26852 21420
rect 27020 21140 27076 21868
rect 27244 21476 27300 21486
rect 27244 21382 27300 21420
rect 27020 21084 27412 21140
rect 27244 20802 27300 20814
rect 27244 20750 27246 20802
rect 27298 20750 27300 20802
rect 26796 20690 26852 20702
rect 26796 20638 26798 20690
rect 26850 20638 26852 20690
rect 26796 20468 26852 20638
rect 27020 20692 27076 20702
rect 27244 20692 27300 20750
rect 27020 20690 27188 20692
rect 27020 20638 27022 20690
rect 27074 20638 27188 20690
rect 27020 20636 27188 20638
rect 27020 20626 27076 20636
rect 26796 20402 26852 20412
rect 26348 20300 26740 20356
rect 26684 20244 26740 20300
rect 26684 20188 26852 20244
rect 26236 20132 26292 20142
rect 26236 20018 26292 20076
rect 26572 20130 26628 20142
rect 26572 20078 26574 20130
rect 26626 20078 26628 20130
rect 26572 20020 26628 20078
rect 26236 19966 26238 20018
rect 26290 19966 26292 20018
rect 26236 19954 26292 19966
rect 26348 19964 26628 20020
rect 26236 19796 26292 19806
rect 26236 19236 26292 19740
rect 26236 19142 26292 19180
rect 26236 17780 26292 17790
rect 26236 17220 26292 17724
rect 26236 17154 26292 17164
rect 26236 16996 26292 17006
rect 26236 14644 26292 16940
rect 26348 15202 26404 19964
rect 26460 19572 26516 19582
rect 26460 16660 26516 19516
rect 26684 19572 26740 19582
rect 26684 18674 26740 19516
rect 26796 19012 26852 20188
rect 27132 19348 27188 20636
rect 27244 20626 27300 20636
rect 27132 19282 27188 19292
rect 27132 19012 27188 19022
rect 26796 19010 27188 19012
rect 26796 18958 27134 19010
rect 27186 18958 27188 19010
rect 26796 18956 27188 18958
rect 26684 18622 26686 18674
rect 26738 18622 26740 18674
rect 26684 18610 26740 18622
rect 26908 17668 26964 17678
rect 26908 17574 26964 17612
rect 26572 17556 26628 17566
rect 26572 16884 26628 17500
rect 26908 17444 26964 17454
rect 26572 16882 26740 16884
rect 26572 16830 26574 16882
rect 26626 16830 26740 16882
rect 26572 16828 26740 16830
rect 26572 16818 26628 16828
rect 26460 16604 26628 16660
rect 26572 15316 26628 16604
rect 26572 15250 26628 15260
rect 26684 16100 26740 16828
rect 26796 16660 26852 16670
rect 26796 16566 26852 16604
rect 26348 15150 26350 15202
rect 26402 15150 26404 15202
rect 26348 15138 26404 15150
rect 26460 15204 26516 15214
rect 26236 14588 26404 14644
rect 26236 14420 26292 14430
rect 26124 14364 26236 14420
rect 26236 14326 26292 14364
rect 26348 13972 26404 14588
rect 25900 13918 25902 13970
rect 25954 13918 25956 13970
rect 25900 13906 25956 13918
rect 26236 13916 26404 13972
rect 26012 13636 26068 13646
rect 25788 11778 25844 11788
rect 25900 13634 26068 13636
rect 25900 13582 26014 13634
rect 26066 13582 26068 13634
rect 25900 13580 26068 13582
rect 25900 11620 25956 13580
rect 26012 13570 26068 13580
rect 26124 12292 26180 12302
rect 26124 12198 26180 12236
rect 25676 11508 25732 11546
rect 25676 11442 25732 11452
rect 25788 11172 25844 11182
rect 25788 11078 25844 11116
rect 25788 10724 25844 10734
rect 25900 10724 25956 11564
rect 25844 10668 25956 10724
rect 26012 12178 26068 12190
rect 26012 12126 26014 12178
rect 26066 12126 26068 12178
rect 25788 10630 25844 10668
rect 25676 10612 25732 10622
rect 25676 9828 25732 10556
rect 26012 10612 26068 12126
rect 26012 10546 26068 10556
rect 26124 11282 26180 11294
rect 26124 11230 26126 11282
rect 26178 11230 26180 11282
rect 26124 10164 26180 11230
rect 26236 10500 26292 13916
rect 26348 13636 26404 13646
rect 26348 12402 26404 13580
rect 26348 12350 26350 12402
rect 26402 12350 26404 12402
rect 26348 12338 26404 12350
rect 26460 12962 26516 15148
rect 26572 14530 26628 14542
rect 26572 14478 26574 14530
rect 26626 14478 26628 14530
rect 26572 14196 26628 14478
rect 26572 14130 26628 14140
rect 26684 13188 26740 16044
rect 26796 16324 26852 16334
rect 26796 16098 26852 16268
rect 26908 16210 26964 17388
rect 27020 16660 27076 18956
rect 27132 18946 27188 18956
rect 27132 18788 27188 18798
rect 27132 18450 27188 18732
rect 27132 18398 27134 18450
rect 27186 18398 27188 18450
rect 27132 18386 27188 18398
rect 27244 17666 27300 17678
rect 27244 17614 27246 17666
rect 27298 17614 27300 17666
rect 27244 17108 27300 17614
rect 27244 17042 27300 17052
rect 27132 16884 27188 16894
rect 27132 16790 27188 16828
rect 27020 16604 27188 16660
rect 26908 16158 26910 16210
rect 26962 16158 26964 16210
rect 26908 16146 26964 16158
rect 26796 16046 26798 16098
rect 26850 16046 26852 16098
rect 26796 16034 26852 16046
rect 27020 15986 27076 15998
rect 27020 15934 27022 15986
rect 27074 15934 27076 15986
rect 26908 15428 26964 15438
rect 26908 14644 26964 15372
rect 26908 14418 26964 14588
rect 26908 14366 26910 14418
rect 26962 14366 26964 14418
rect 26908 14354 26964 14366
rect 27020 13746 27076 15934
rect 27132 15876 27188 16604
rect 27132 15810 27188 15820
rect 27132 14420 27188 14430
rect 27132 14326 27188 14364
rect 27020 13694 27022 13746
rect 27074 13694 27076 13746
rect 27020 13682 27076 13694
rect 27132 13858 27188 13870
rect 27132 13806 27134 13858
rect 27186 13806 27188 13858
rect 26908 13300 26964 13310
rect 26684 13132 26852 13188
rect 26684 12964 26740 12974
rect 26460 12910 26462 12962
rect 26514 12910 26516 12962
rect 26460 11620 26516 12910
rect 26572 12962 26740 12964
rect 26572 12910 26686 12962
rect 26738 12910 26740 12962
rect 26572 12908 26740 12910
rect 26572 11844 26628 12908
rect 26684 12898 26740 12908
rect 26572 11778 26628 11788
rect 26684 12404 26740 12414
rect 26796 12404 26852 13132
rect 26684 12402 26852 12404
rect 26684 12350 26686 12402
rect 26738 12350 26852 12402
rect 26684 12348 26852 12350
rect 26348 11564 26516 11620
rect 26348 10724 26404 11564
rect 26460 11394 26516 11406
rect 26460 11342 26462 11394
rect 26514 11342 26516 11394
rect 26460 11282 26516 11342
rect 26460 11230 26462 11282
rect 26514 11230 26516 11282
rect 26460 11218 26516 11230
rect 26572 11396 26628 11406
rect 26572 11170 26628 11340
rect 26572 11118 26574 11170
rect 26626 11118 26628 11170
rect 26572 11106 26628 11118
rect 26348 10668 26516 10724
rect 26348 10500 26404 10510
rect 26236 10498 26404 10500
rect 26236 10446 26350 10498
rect 26402 10446 26404 10498
rect 26236 10444 26404 10446
rect 26348 10386 26404 10444
rect 26348 10334 26350 10386
rect 26402 10334 26404 10386
rect 26348 10322 26404 10334
rect 26460 10276 26516 10668
rect 26460 10220 26628 10276
rect 26124 10108 26516 10164
rect 25788 10052 25844 10062
rect 25788 10050 26068 10052
rect 25788 9998 25790 10050
rect 25842 9998 26068 10050
rect 25788 9996 26068 9998
rect 25788 9986 25844 9996
rect 25676 9772 25956 9828
rect 25340 8642 25396 8652
rect 25452 9548 25620 9604
rect 25676 9602 25732 9614
rect 25676 9550 25678 9602
rect 25730 9550 25732 9602
rect 25228 8306 25284 8316
rect 25340 7588 25396 7598
rect 25340 7494 25396 7532
rect 25340 7028 25396 7038
rect 25340 6690 25396 6972
rect 25340 6638 25342 6690
rect 25394 6638 25396 6690
rect 25340 6626 25396 6638
rect 25340 6244 25396 6254
rect 25340 6130 25396 6188
rect 25340 6078 25342 6130
rect 25394 6078 25396 6130
rect 25340 6066 25396 6078
rect 25452 6130 25508 9548
rect 25676 9380 25732 9550
rect 25788 9380 25844 9390
rect 25564 9324 25788 9380
rect 25564 9042 25620 9324
rect 25788 9314 25844 9324
rect 25564 8990 25566 9042
rect 25618 8990 25620 9042
rect 25564 8978 25620 8990
rect 25676 9044 25732 9054
rect 25676 8950 25732 8988
rect 25900 9042 25956 9772
rect 25900 8990 25902 9042
rect 25954 8990 25956 9042
rect 25788 8930 25844 8942
rect 25788 8878 25790 8930
rect 25842 8878 25844 8930
rect 25788 8596 25844 8878
rect 25788 8530 25844 8540
rect 25900 8372 25956 8990
rect 26012 9266 26068 9996
rect 26460 10050 26516 10108
rect 26460 9998 26462 10050
rect 26514 9998 26516 10050
rect 26460 9986 26516 9998
rect 26460 9826 26516 9838
rect 26460 9774 26462 9826
rect 26514 9774 26516 9826
rect 26012 9214 26014 9266
rect 26066 9214 26068 9266
rect 26012 8932 26068 9214
rect 26124 9714 26180 9726
rect 26124 9662 26126 9714
rect 26178 9662 26180 9714
rect 26124 9268 26180 9662
rect 26460 9380 26516 9774
rect 26572 9716 26628 10220
rect 26572 9650 26628 9660
rect 26460 9314 26516 9324
rect 26124 9202 26180 9212
rect 26572 9156 26628 9166
rect 26460 9042 26516 9054
rect 26460 8990 26462 9042
rect 26514 8990 26516 9042
rect 26460 8932 26516 8990
rect 26012 8876 26516 8932
rect 25788 8316 25956 8372
rect 26012 8708 26068 8718
rect 25788 8148 25844 8316
rect 25788 8082 25844 8092
rect 25900 8036 25956 8046
rect 26012 8036 26068 8652
rect 25900 8034 26068 8036
rect 25900 7982 25902 8034
rect 25954 7982 26068 8034
rect 25900 7980 26068 7982
rect 26348 8036 26404 8046
rect 25900 7970 25956 7980
rect 26348 7942 26404 7980
rect 26012 7588 26068 7598
rect 26012 7494 26068 7532
rect 25676 7474 25732 7486
rect 25676 7422 25678 7474
rect 25730 7422 25732 7474
rect 25676 7028 25732 7422
rect 26236 7476 26292 7486
rect 26012 7364 26068 7374
rect 26012 7270 26068 7308
rect 25676 6962 25732 6972
rect 25900 7140 25956 7150
rect 25452 6078 25454 6130
rect 25506 6078 25508 6130
rect 25004 5628 25172 5684
rect 25228 5906 25284 5918
rect 25228 5854 25230 5906
rect 25282 5854 25284 5906
rect 24108 5394 24164 5404
rect 24780 5572 24836 5582
rect 23884 5182 23886 5234
rect 23938 5182 23940 5234
rect 23884 5170 23940 5182
rect 24332 5348 24388 5358
rect 24332 5234 24388 5292
rect 24332 5182 24334 5234
rect 24386 5182 24388 5234
rect 24332 5170 24388 5182
rect 24780 5122 24836 5516
rect 24780 5070 24782 5122
rect 24834 5070 24836 5122
rect 24332 4564 24388 4574
rect 23772 4562 24332 4564
rect 23772 4510 23774 4562
rect 23826 4510 24332 4562
rect 23772 4508 24332 4510
rect 23772 4498 23828 4508
rect 24332 4470 24388 4508
rect 24668 4564 24724 4574
rect 24780 4564 24836 5070
rect 24668 4562 24836 4564
rect 24668 4510 24670 4562
rect 24722 4510 24836 4562
rect 24668 4508 24836 4510
rect 24668 4498 24724 4508
rect 23436 4452 23492 4462
rect 23324 4450 23492 4452
rect 23324 4398 23438 4450
rect 23490 4398 23492 4450
rect 23324 4396 23492 4398
rect 22876 4386 22932 4396
rect 22764 4286 22766 4338
rect 22818 4286 22820 4338
rect 22764 4274 22820 4286
rect 22988 4116 23044 4126
rect 23100 4116 23156 4126
rect 22988 4114 23100 4116
rect 22988 4062 22990 4114
rect 23042 4062 23100 4114
rect 22988 4060 23100 4062
rect 22988 4050 23044 4060
rect 22540 3836 23044 3892
rect 20972 3614 20974 3666
rect 21026 3614 21028 3666
rect 20188 3602 20244 3612
rect 20972 3602 21028 3614
rect 21308 3778 21364 3790
rect 21308 3726 21310 3778
rect 21362 3726 21364 3778
rect 21308 3666 21364 3726
rect 21308 3614 21310 3666
rect 21362 3614 21364 3666
rect 21308 3602 21364 3614
rect 22988 3666 23044 3836
rect 22988 3614 22990 3666
rect 23042 3614 23044 3666
rect 22988 3602 23044 3614
rect 21980 3556 22036 3566
rect 21980 3462 22036 3500
rect 23100 3556 23156 4060
rect 23436 3666 23492 4396
rect 23436 3614 23438 3666
rect 23490 3614 23492 3666
rect 23436 3602 23492 3614
rect 23100 3490 23156 3500
rect 19740 3266 19796 3276
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 25004 2884 25060 5628
rect 25228 5348 25284 5854
rect 25452 5348 25508 6078
rect 25228 5282 25284 5292
rect 25340 5292 25452 5348
rect 25116 5234 25172 5246
rect 25116 5182 25118 5234
rect 25170 5182 25172 5234
rect 25116 5124 25172 5182
rect 25116 5058 25172 5068
rect 25340 4676 25396 5292
rect 25452 5282 25508 5292
rect 25564 6466 25620 6478
rect 25564 6414 25566 6466
rect 25618 6414 25620 6466
rect 25452 5122 25508 5134
rect 25452 5070 25454 5122
rect 25506 5070 25508 5122
rect 25452 5012 25508 5070
rect 25452 4946 25508 4956
rect 25340 4610 25396 4620
rect 25452 4564 25508 4574
rect 25452 4470 25508 4508
rect 25228 4452 25284 4462
rect 25228 4358 25284 4396
rect 25564 4452 25620 6414
rect 25788 6356 25844 6366
rect 25788 5572 25844 6300
rect 25900 5908 25956 7084
rect 26236 6580 26292 7420
rect 26572 6916 26628 9100
rect 26684 8820 26740 12348
rect 26908 11956 26964 13244
rect 26908 10724 26964 11900
rect 26796 10668 26964 10724
rect 27020 11060 27076 11070
rect 26796 9716 26852 10668
rect 27020 10610 27076 11004
rect 27132 10722 27188 13806
rect 27244 13188 27300 13198
rect 27244 13074 27300 13132
rect 27244 13022 27246 13074
rect 27298 13022 27300 13074
rect 27244 13010 27300 13022
rect 27356 12740 27412 21084
rect 27468 20132 27524 21868
rect 27692 20692 27748 22092
rect 27804 21810 27860 22092
rect 27916 22036 27972 25340
rect 28028 22932 28084 26572
rect 28252 26290 28308 26302
rect 28252 26238 28254 26290
rect 28306 26238 28308 26290
rect 28140 25956 28196 25966
rect 28140 25618 28196 25900
rect 28140 25566 28142 25618
rect 28194 25566 28196 25618
rect 28140 25554 28196 25566
rect 28252 25508 28308 26238
rect 28476 26068 28532 26078
rect 28476 25974 28532 26012
rect 28252 25172 28308 25452
rect 28588 25508 28644 26796
rect 28924 26404 28980 27580
rect 29148 27076 29204 27086
rect 29148 26982 29204 27020
rect 29260 26964 29316 28028
rect 29876 28028 30212 28084
rect 29820 27990 29876 28028
rect 29260 26898 29316 26908
rect 29372 27186 29428 27198
rect 29372 27134 29374 27186
rect 29426 27134 29428 27186
rect 28924 26348 29204 26404
rect 29148 26290 29204 26348
rect 29148 26238 29150 26290
rect 29202 26238 29204 26290
rect 29148 25844 29204 26238
rect 29148 25778 29204 25788
rect 29372 26292 29428 27134
rect 30156 27074 30212 28028
rect 30828 28082 30940 28084
rect 30828 28030 30830 28082
rect 30882 28030 30940 28082
rect 30828 28028 30940 28030
rect 30828 28018 30884 28028
rect 30940 27990 30996 28028
rect 31276 28420 31332 28430
rect 30156 27022 30158 27074
rect 30210 27022 30212 27074
rect 30156 27010 30212 27022
rect 31276 27074 31332 28364
rect 32396 28308 32452 35084
rect 33292 35074 33348 35084
rect 33516 35028 33572 35038
rect 33628 35028 33684 35646
rect 34076 35140 34132 35150
rect 33852 35028 33908 35038
rect 33572 35026 33908 35028
rect 33572 34974 33854 35026
rect 33906 34974 33908 35026
rect 33572 34972 33908 34974
rect 33516 34962 33572 34972
rect 33852 34962 33908 34972
rect 32732 34804 32788 34814
rect 32732 34710 32788 34748
rect 33516 34802 33572 34814
rect 33516 34750 33518 34802
rect 33570 34750 33572 34802
rect 32844 34690 32900 34702
rect 32844 34638 32846 34690
rect 32898 34638 32900 34690
rect 32844 34132 32900 34638
rect 33516 34356 33572 34750
rect 34076 34580 34132 35084
rect 34188 35028 34244 36206
rect 34524 35924 34580 36764
rect 34860 36708 34916 36718
rect 34860 35924 34916 36652
rect 34412 35868 34580 35924
rect 34636 35868 34860 35924
rect 34300 35476 34356 35486
rect 34300 35382 34356 35420
rect 34412 35364 34468 35868
rect 34524 35700 34580 35710
rect 34524 35606 34580 35644
rect 34412 35298 34468 35308
rect 34188 34972 34468 35028
rect 34188 34692 34244 34702
rect 34188 34690 34356 34692
rect 34188 34638 34190 34690
rect 34242 34638 34356 34690
rect 34188 34636 34356 34638
rect 34188 34626 34244 34636
rect 34076 34514 34132 34524
rect 33516 34290 33572 34300
rect 34188 34356 34244 34366
rect 34188 34262 34244 34300
rect 33628 34244 33684 34254
rect 33628 34150 33684 34188
rect 32844 34066 32900 34076
rect 34300 33348 34356 34636
rect 34412 34132 34468 34972
rect 34412 34066 34468 34076
rect 34636 33572 34692 35868
rect 34860 35830 34916 35868
rect 34972 34356 35028 37886
rect 35532 37604 35588 38782
rect 36092 38834 36148 38846
rect 36092 38782 36094 38834
rect 36146 38782 36148 38834
rect 35644 38724 35700 38734
rect 35644 37938 35700 38668
rect 35980 38722 36036 38734
rect 35980 38670 35982 38722
rect 36034 38670 36036 38722
rect 35644 37886 35646 37938
rect 35698 37886 35700 37938
rect 35644 37874 35700 37886
rect 35756 38162 35812 38174
rect 35756 38110 35758 38162
rect 35810 38110 35812 38162
rect 35756 37828 35812 38110
rect 35756 37762 35812 37772
rect 35868 38050 35924 38062
rect 35868 37998 35870 38050
rect 35922 37998 35924 38050
rect 35532 37538 35588 37548
rect 35644 37492 35700 37502
rect 35084 37380 35140 37390
rect 35084 36706 35140 37324
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35084 36654 35086 36706
rect 35138 36654 35140 36706
rect 35084 36642 35140 36654
rect 35420 36708 35476 36718
rect 35420 36614 35476 36652
rect 35196 36482 35252 36494
rect 35196 36430 35198 36482
rect 35250 36430 35252 36482
rect 35196 36148 35252 36430
rect 35196 36082 35252 36092
rect 35644 36482 35700 37436
rect 35644 36430 35646 36482
rect 35698 36430 35700 36482
rect 35308 35700 35364 35710
rect 35644 35700 35700 36430
rect 35868 35812 35924 37998
rect 35980 37716 36036 38670
rect 36092 37940 36148 38782
rect 36316 38668 36372 39004
rect 36092 37874 36148 37884
rect 36204 38612 36372 38668
rect 35980 37650 36036 37660
rect 36204 37266 36260 38612
rect 36204 37214 36206 37266
rect 36258 37214 36260 37266
rect 36204 37202 36260 37214
rect 36092 36708 36148 36718
rect 36092 36614 36148 36652
rect 36428 36484 36484 39676
rect 36092 36428 36484 36484
rect 35980 36372 36036 36382
rect 35980 36278 36036 36316
rect 36092 36370 36148 36428
rect 36092 36318 36094 36370
rect 36146 36318 36148 36370
rect 35308 35698 35700 35700
rect 35308 35646 35310 35698
rect 35362 35646 35700 35698
rect 35308 35644 35700 35646
rect 35756 35700 35812 35710
rect 35868 35700 35924 35756
rect 35756 35698 35924 35700
rect 35756 35646 35758 35698
rect 35810 35646 35924 35698
rect 35756 35644 35924 35646
rect 36092 35700 36148 36318
rect 35308 35634 35364 35644
rect 35756 35634 35812 35644
rect 36092 35634 36148 35644
rect 36204 35924 36260 35934
rect 36204 35810 36260 35868
rect 36204 35758 36206 35810
rect 36258 35758 36260 35810
rect 35756 35364 35812 35374
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 34972 34290 35028 34300
rect 35756 34354 35812 35308
rect 35756 34302 35758 34354
rect 35810 34302 35812 34354
rect 35756 34290 35812 34302
rect 34860 34244 34916 34254
rect 34860 34150 34916 34188
rect 34748 34132 34804 34142
rect 36204 34132 36260 35758
rect 36316 35474 36372 35486
rect 36316 35422 36318 35474
rect 36370 35422 36372 35474
rect 36316 34916 36372 35422
rect 36316 34850 36372 34860
rect 36316 34132 36372 34142
rect 36204 34130 36372 34132
rect 36204 34078 36318 34130
rect 36370 34078 36372 34130
rect 36204 34076 36372 34078
rect 34748 34038 34804 34076
rect 36316 34066 36372 34076
rect 36428 33908 36484 33918
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 34300 33282 34356 33292
rect 34412 33516 34692 33572
rect 34300 33124 34356 33134
rect 34412 33124 34468 33516
rect 34300 33122 34468 33124
rect 34300 33070 34302 33122
rect 34354 33070 34468 33122
rect 34300 33068 34468 33070
rect 36204 33346 36260 33358
rect 36204 33294 36206 33346
rect 36258 33294 36260 33346
rect 34300 33058 34356 33068
rect 36204 32788 36260 33294
rect 36428 33234 36484 33852
rect 36428 33182 36430 33234
rect 36482 33182 36484 33234
rect 36428 33170 36484 33182
rect 36204 32722 36260 32732
rect 33628 32562 33684 32574
rect 33628 32510 33630 32562
rect 33682 32510 33684 32562
rect 32732 32004 32788 32014
rect 32732 31666 32788 31948
rect 32732 31614 32734 31666
rect 32786 31614 32788 31666
rect 32732 31602 32788 31614
rect 32956 31668 33012 31678
rect 32956 31108 33012 31612
rect 33516 31556 33572 31566
rect 32956 31042 33012 31052
rect 33068 31554 33572 31556
rect 33068 31502 33518 31554
rect 33570 31502 33572 31554
rect 33068 31500 33572 31502
rect 32396 28242 32452 28252
rect 32620 30212 32676 30222
rect 32620 28082 32676 30156
rect 32732 30210 32788 30222
rect 32732 30158 32734 30210
rect 32786 30158 32788 30210
rect 32732 30100 32788 30158
rect 32732 30034 32788 30044
rect 32844 30100 32900 30110
rect 33068 30100 33124 31500
rect 32844 30098 33124 30100
rect 32844 30046 32846 30098
rect 32898 30046 33124 30098
rect 32844 30044 33124 30046
rect 33180 31332 33236 31342
rect 32844 30034 32900 30044
rect 33068 29428 33124 29438
rect 33068 28754 33124 29372
rect 33180 29426 33236 31276
rect 33516 30994 33572 31500
rect 33628 31332 33684 32510
rect 34076 32562 34132 32574
rect 34076 32510 34078 32562
rect 34130 32510 34132 32562
rect 33740 31778 33796 31790
rect 33740 31726 33742 31778
rect 33794 31726 33796 31778
rect 33740 31668 33796 31726
rect 33740 31602 33796 31612
rect 34076 31554 34132 32510
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 34188 31780 34244 31790
rect 34188 31686 34244 31724
rect 34300 31778 34356 31790
rect 34300 31726 34302 31778
rect 34354 31726 34356 31778
rect 34076 31502 34078 31554
rect 34130 31502 34132 31554
rect 34076 31490 34132 31502
rect 34300 31332 34356 31726
rect 33628 31266 33684 31276
rect 33740 31276 34356 31332
rect 33740 31218 33796 31276
rect 33740 31166 33742 31218
rect 33794 31166 33796 31218
rect 33740 31154 33796 31166
rect 36540 31220 36596 40908
rect 36652 35140 36708 42252
rect 36876 38668 36932 45500
rect 36988 43540 37044 46508
rect 37100 44436 37156 46956
rect 37100 44370 37156 44380
rect 37324 43652 37380 48412
rect 37548 48356 37604 48974
rect 37884 48916 37940 48926
rect 37884 48822 37940 48860
rect 37772 48356 37828 48366
rect 37996 48356 38052 49084
rect 38108 48468 38164 49644
rect 38444 49140 38500 49980
rect 38444 49026 38500 49084
rect 38444 48974 38446 49026
rect 38498 48974 38500 49026
rect 38444 48962 38500 48974
rect 38332 48916 38388 48926
rect 38332 48822 38388 48860
rect 38556 48914 38612 48926
rect 38556 48862 38558 48914
rect 38610 48862 38612 48914
rect 38220 48468 38276 48478
rect 38108 48412 38220 48468
rect 37548 48354 37828 48356
rect 37548 48302 37774 48354
rect 37826 48302 37828 48354
rect 37548 48300 37828 48302
rect 37436 47460 37492 47470
rect 37436 47366 37492 47404
rect 37548 47236 37604 48300
rect 37772 48290 37828 48300
rect 37884 48354 38052 48356
rect 37884 48302 37998 48354
rect 38050 48302 38052 48354
rect 37884 48300 38052 48302
rect 37660 48132 37716 48142
rect 37660 48038 37716 48076
rect 37884 47908 37940 48300
rect 37996 48290 38052 48300
rect 38220 48242 38276 48412
rect 38556 48468 38612 48862
rect 38556 48402 38612 48412
rect 38220 48190 38222 48242
rect 38274 48190 38276 48242
rect 37660 47852 37940 47908
rect 38108 48020 38164 48030
rect 37660 47458 37716 47852
rect 37660 47406 37662 47458
rect 37714 47406 37716 47458
rect 37660 47394 37716 47406
rect 38108 47458 38164 47964
rect 38108 47406 38110 47458
rect 38162 47406 38164 47458
rect 38108 47394 38164 47406
rect 38220 47460 38276 48190
rect 38668 48020 38724 48030
rect 38668 47926 38724 47964
rect 38220 47394 38276 47404
rect 37884 47236 37940 47246
rect 37548 47234 37940 47236
rect 37548 47182 37886 47234
rect 37938 47182 37940 47234
rect 37548 47180 37940 47182
rect 37884 46340 37940 47180
rect 38220 47236 38276 47246
rect 38220 47234 38612 47236
rect 38220 47182 38222 47234
rect 38274 47182 38612 47234
rect 38220 47180 38612 47182
rect 38220 47170 38276 47180
rect 38444 47012 38500 47022
rect 37996 46564 38052 46574
rect 37996 46470 38052 46508
rect 38444 46564 38500 46956
rect 38444 46470 38500 46508
rect 37660 46284 37940 46340
rect 37548 44322 37604 44334
rect 37548 44270 37550 44322
rect 37602 44270 37604 44322
rect 37548 44212 37604 44270
rect 37548 44146 37604 44156
rect 37436 43652 37492 43662
rect 37324 43596 37436 43652
rect 37436 43586 37492 43596
rect 37548 43540 37604 43550
rect 36988 43484 37156 43540
rect 36988 41074 37044 41086
rect 36988 41022 36990 41074
rect 37042 41022 37044 41074
rect 36988 40628 37044 41022
rect 36988 40562 37044 40572
rect 37100 38668 37156 43484
rect 37212 43316 37268 43326
rect 37212 43314 37380 43316
rect 37212 43262 37214 43314
rect 37266 43262 37380 43314
rect 37212 43260 37380 43262
rect 37212 43250 37268 43260
rect 37212 41186 37268 41198
rect 37212 41134 37214 41186
rect 37266 41134 37268 41186
rect 37212 40964 37268 41134
rect 37212 40898 37268 40908
rect 37324 39842 37380 43260
rect 37324 39790 37326 39842
rect 37378 39790 37380 39842
rect 37324 39778 37380 39790
rect 37436 42754 37492 42766
rect 37436 42702 37438 42754
rect 37490 42702 37492 42754
rect 37436 39620 37492 42702
rect 37548 42754 37604 43484
rect 37548 42702 37550 42754
rect 37602 42702 37604 42754
rect 37548 42690 37604 42702
rect 37548 41412 37604 41422
rect 37660 41412 37716 46284
rect 38556 45890 38612 47180
rect 38780 47012 38836 47022
rect 38780 46898 38836 46956
rect 38780 46846 38782 46898
rect 38834 46846 38836 46898
rect 38780 46834 38836 46846
rect 38556 45838 38558 45890
rect 38610 45838 38612 45890
rect 38556 45826 38612 45838
rect 38780 45668 38836 45678
rect 38780 45574 38836 45612
rect 38892 45444 38948 50372
rect 39340 49812 39396 49822
rect 39004 49810 39396 49812
rect 39004 49758 39342 49810
rect 39394 49758 39396 49810
rect 39004 49756 39396 49758
rect 39004 49250 39060 49756
rect 39340 49746 39396 49756
rect 39004 49198 39006 49250
rect 39058 49198 39060 49250
rect 39004 49186 39060 49198
rect 39452 49028 39508 50372
rect 39340 49026 39508 49028
rect 39340 48974 39454 49026
rect 39506 48974 39508 49026
rect 39340 48972 39508 48974
rect 39004 48468 39060 48478
rect 39004 48374 39060 48412
rect 39340 47572 39396 48972
rect 39452 48962 39508 48972
rect 39564 49028 39620 50652
rect 39676 50706 39732 51212
rect 40236 51154 40292 52108
rect 40236 51102 40238 51154
rect 40290 51102 40292 51154
rect 40236 51090 40292 51102
rect 40348 51378 40404 51390
rect 40348 51326 40350 51378
rect 40402 51326 40404 51378
rect 39676 50654 39678 50706
rect 39730 50654 39732 50706
rect 39676 50642 39732 50654
rect 40236 49812 40292 49822
rect 40236 49718 40292 49756
rect 39788 49698 39844 49710
rect 39788 49646 39790 49698
rect 39842 49646 39844 49698
rect 39788 49138 39844 49646
rect 40348 49252 40404 51326
rect 40460 50260 40516 57148
rect 40460 50194 40516 50204
rect 40572 50036 40628 57372
rect 41020 55970 41076 59200
rect 45724 56308 45780 59200
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 45724 56242 45780 56252
rect 48412 56308 48468 56318
rect 48412 56214 48468 56252
rect 41020 55918 41022 55970
rect 41074 55918 41076 55970
rect 41020 55906 41076 55918
rect 41692 56084 41748 56094
rect 40908 55298 40964 55310
rect 40908 55246 40910 55298
rect 40962 55246 40964 55298
rect 40908 54628 40964 55246
rect 41020 55188 41076 55198
rect 41356 55188 41412 55198
rect 41020 55186 41412 55188
rect 41020 55134 41022 55186
rect 41074 55134 41358 55186
rect 41410 55134 41412 55186
rect 41020 55132 41412 55134
rect 41020 55122 41076 55132
rect 41356 55122 41412 55132
rect 41692 55186 41748 56028
rect 42588 56084 42644 56094
rect 42588 55990 42644 56028
rect 46508 56084 46564 56094
rect 41692 55134 41694 55186
rect 41746 55134 41748 55186
rect 41692 55122 41748 55134
rect 41804 55300 41860 55310
rect 40908 54572 41300 54628
rect 41244 54516 41300 54572
rect 41244 54514 41524 54516
rect 41244 54462 41246 54514
rect 41298 54462 41524 54514
rect 41244 54460 41524 54462
rect 41244 54450 41300 54460
rect 40684 53956 40740 53966
rect 40684 53862 40740 53900
rect 41468 53954 41524 54460
rect 41804 54514 41860 55244
rect 43372 55300 43428 55310
rect 43372 55206 43428 55244
rect 43820 55298 43876 55310
rect 43820 55246 43822 55298
rect 43874 55246 43876 55298
rect 42476 55188 42532 55198
rect 42476 55094 42532 55132
rect 42700 55188 42756 55198
rect 42700 55094 42756 55132
rect 43820 55188 43876 55246
rect 44044 55300 44100 55310
rect 44940 55300 44996 55310
rect 44044 55298 45108 55300
rect 44044 55246 44046 55298
rect 44098 55246 44942 55298
rect 44994 55246 45108 55298
rect 44044 55244 45108 55246
rect 44044 55234 44100 55244
rect 44940 55234 44996 55244
rect 42252 55076 42308 55086
rect 42588 55076 42644 55086
rect 42252 55074 42420 55076
rect 42252 55022 42254 55074
rect 42306 55022 42420 55074
rect 42252 55020 42420 55022
rect 42252 55010 42308 55020
rect 42364 54740 42420 55020
rect 42588 54982 42644 55020
rect 42364 54684 43428 54740
rect 41804 54462 41806 54514
rect 41858 54462 41860 54514
rect 41804 54450 41860 54462
rect 42028 54514 42084 54526
rect 42028 54462 42030 54514
rect 42082 54462 42084 54514
rect 41916 54402 41972 54414
rect 41916 54350 41918 54402
rect 41970 54350 41972 54402
rect 41916 54292 41972 54350
rect 41916 54226 41972 54236
rect 41468 53902 41470 53954
rect 41522 53902 41524 53954
rect 41468 53890 41524 53902
rect 42028 53956 42084 54462
rect 42140 54516 42196 54526
rect 42140 54422 42196 54460
rect 42700 54514 42756 54526
rect 42700 54462 42702 54514
rect 42754 54462 42756 54514
rect 42700 54404 42756 54462
rect 42700 54338 42756 54348
rect 42812 54516 42868 54526
rect 42028 53890 42084 53900
rect 42812 53954 42868 54460
rect 42812 53902 42814 53954
rect 42866 53902 42868 53954
rect 42812 53890 42868 53902
rect 43260 53954 43316 54684
rect 43372 54514 43428 54684
rect 43372 54462 43374 54514
rect 43426 54462 43428 54514
rect 43372 54450 43428 54462
rect 43708 54516 43764 54526
rect 43708 54422 43764 54460
rect 43820 54402 43876 55132
rect 43820 54350 43822 54402
rect 43874 54350 43876 54402
rect 43820 54338 43876 54350
rect 43932 54626 43988 54638
rect 43932 54574 43934 54626
rect 43986 54574 43988 54626
rect 43260 53902 43262 53954
rect 43314 53902 43316 53954
rect 43260 53890 43316 53902
rect 40796 53844 40852 53854
rect 40796 53750 40852 53788
rect 42252 53732 42308 53742
rect 42252 53638 42308 53676
rect 42476 53730 42532 53742
rect 42476 53678 42478 53730
rect 42530 53678 42532 53730
rect 41356 53620 41412 53630
rect 41356 53526 41412 53564
rect 42476 53620 42532 53678
rect 43260 53732 43316 53742
rect 40908 53506 40964 53518
rect 40908 53454 40910 53506
rect 40962 53454 40964 53506
rect 40908 51604 40964 53454
rect 41468 53506 41524 53518
rect 41468 53454 41470 53506
rect 41522 53454 41524 53506
rect 41468 52836 41524 53454
rect 41804 52836 41860 52846
rect 41468 52834 41860 52836
rect 41468 52782 41806 52834
rect 41858 52782 41860 52834
rect 41468 52780 41860 52782
rect 41244 52388 41300 52398
rect 41020 52276 41076 52286
rect 41020 52162 41076 52220
rect 41020 52110 41022 52162
rect 41074 52110 41076 52162
rect 41020 52098 41076 52110
rect 41132 52164 41188 52174
rect 41132 52070 41188 52108
rect 41244 52162 41300 52332
rect 41692 52388 41748 52398
rect 41692 52294 41748 52332
rect 41244 52110 41246 52162
rect 41298 52110 41300 52162
rect 41244 52098 41300 52110
rect 40908 51538 40964 51548
rect 41692 51268 41748 51278
rect 40572 49970 40628 49980
rect 41020 50260 41076 50270
rect 41020 50034 41076 50204
rect 41020 49982 41022 50034
rect 41074 49982 41076 50034
rect 41020 49970 41076 49982
rect 41468 50036 41524 50046
rect 41468 49942 41524 49980
rect 40348 49186 40404 49196
rect 39788 49086 39790 49138
rect 39842 49086 39844 49138
rect 39788 49074 39844 49086
rect 41692 49138 41748 51212
rect 41692 49086 41694 49138
rect 41746 49086 41748 49138
rect 41692 49074 41748 49086
rect 40796 49028 40852 49038
rect 39564 48934 39620 48972
rect 40124 49026 40852 49028
rect 40124 48974 40798 49026
rect 40850 48974 40852 49026
rect 40124 48972 40852 48974
rect 39900 48916 39956 48926
rect 39900 48242 39956 48860
rect 40124 48466 40180 48972
rect 40796 48962 40852 48972
rect 40908 49028 40964 49038
rect 40460 48804 40516 48814
rect 40516 48748 40628 48804
rect 40460 48710 40516 48748
rect 40124 48414 40126 48466
rect 40178 48414 40180 48466
rect 40124 48402 40180 48414
rect 39900 48190 39902 48242
rect 39954 48190 39956 48242
rect 39900 48178 39956 48190
rect 39452 48132 39508 48142
rect 39452 48038 39508 48076
rect 40236 48020 40292 48030
rect 39116 47516 39340 47572
rect 39116 46898 39172 47516
rect 39340 47478 39396 47516
rect 40124 48018 40292 48020
rect 40124 47966 40238 48018
rect 40290 47966 40292 48018
rect 40124 47964 40292 47966
rect 40124 47460 40180 47964
rect 40236 47954 40292 47964
rect 40348 48020 40404 48030
rect 39676 47404 40180 47460
rect 40236 47572 40292 47582
rect 40236 47458 40292 47516
rect 40236 47406 40238 47458
rect 40290 47406 40292 47458
rect 39116 46846 39118 46898
rect 39170 46846 39172 46898
rect 39116 46834 39172 46846
rect 39228 47234 39284 47246
rect 39228 47182 39230 47234
rect 39282 47182 39284 47234
rect 39228 46004 39284 47182
rect 39116 45948 39284 46004
rect 39004 45780 39060 45790
rect 39116 45780 39172 45948
rect 39004 45778 39172 45780
rect 39004 45726 39006 45778
rect 39058 45726 39172 45778
rect 39004 45724 39172 45726
rect 39004 45714 39060 45724
rect 38780 45388 38948 45444
rect 38332 44994 38388 45006
rect 38332 44942 38334 44994
rect 38386 44942 38388 44994
rect 37884 44434 37940 44446
rect 37884 44382 37886 44434
rect 37938 44382 37940 44434
rect 37772 43540 37828 43550
rect 37772 43446 37828 43484
rect 37772 42868 37828 42878
rect 37884 42868 37940 44382
rect 38220 44436 38276 44446
rect 38220 44342 38276 44380
rect 37772 42866 37940 42868
rect 37772 42814 37774 42866
rect 37826 42814 37940 42866
rect 37772 42812 37940 42814
rect 37996 44324 38052 44334
rect 37996 42868 38052 44268
rect 38332 44324 38388 44942
rect 38332 44258 38388 44268
rect 38780 44210 38836 45388
rect 39004 44324 39060 44334
rect 39004 44230 39060 44268
rect 38780 44158 38782 44210
rect 38834 44158 38836 44210
rect 38780 44146 38836 44158
rect 38668 43652 38724 43662
rect 37772 42802 37828 42812
rect 37996 42802 38052 42812
rect 38444 43426 38500 43438
rect 38444 43374 38446 43426
rect 38498 43374 38500 43426
rect 38444 42866 38500 43374
rect 38556 43428 38612 43438
rect 38556 43334 38612 43372
rect 38444 42814 38446 42866
rect 38498 42814 38500 42866
rect 38444 42802 38500 42814
rect 38556 42756 38612 42766
rect 38668 42756 38724 43596
rect 38556 42754 38724 42756
rect 38556 42702 38558 42754
rect 38610 42702 38724 42754
rect 38556 42700 38724 42702
rect 37884 42644 37940 42654
rect 38220 42644 38276 42654
rect 37940 42642 38276 42644
rect 37940 42590 38222 42642
rect 38274 42590 38276 42642
rect 37940 42588 38276 42590
rect 37884 42550 37940 42588
rect 38220 42578 38276 42588
rect 38556 42532 38612 42700
rect 38556 42466 38612 42476
rect 38892 42532 38948 42542
rect 39004 42532 39060 42542
rect 38948 42530 39060 42532
rect 38948 42478 39006 42530
rect 39058 42478 39060 42530
rect 38948 42476 39060 42478
rect 37548 41410 37716 41412
rect 37548 41358 37550 41410
rect 37602 41358 37716 41410
rect 37548 41356 37716 41358
rect 37996 41860 38052 41870
rect 37548 41346 37604 41356
rect 37996 40290 38052 41804
rect 38780 41186 38836 41198
rect 38780 41134 38782 41186
rect 38834 41134 38836 41186
rect 38668 41076 38724 41086
rect 37996 40238 37998 40290
rect 38050 40238 38052 40290
rect 37996 40226 38052 40238
rect 38332 40402 38388 40414
rect 38332 40350 38334 40402
rect 38386 40350 38388 40402
rect 37548 39844 37604 39854
rect 37996 39844 38052 39854
rect 37548 39842 38052 39844
rect 37548 39790 37550 39842
rect 37602 39790 37998 39842
rect 38050 39790 38052 39842
rect 37548 39788 38052 39790
rect 37548 39778 37604 39788
rect 37772 39620 37828 39630
rect 37436 39618 37828 39620
rect 37436 39566 37774 39618
rect 37826 39566 37828 39618
rect 37436 39564 37828 39566
rect 36876 38612 37044 38668
rect 37100 38612 37380 38668
rect 36988 37492 37044 38612
rect 37044 37436 37268 37492
rect 36988 37398 37044 37436
rect 37212 37378 37268 37436
rect 37212 37326 37214 37378
rect 37266 37326 37268 37378
rect 37212 37314 37268 37326
rect 36764 35924 36820 35934
rect 36764 35830 36820 35868
rect 36652 35074 36708 35084
rect 37212 35698 37268 35710
rect 37212 35646 37214 35698
rect 37266 35646 37268 35698
rect 37212 34802 37268 35646
rect 37324 35252 37380 38612
rect 37548 38050 37604 38062
rect 37548 37998 37550 38050
rect 37602 37998 37604 38050
rect 37548 37940 37604 37998
rect 37548 37874 37604 37884
rect 37660 37492 37716 37502
rect 37660 37398 37716 37436
rect 37772 36596 37828 39564
rect 37884 38050 37940 39788
rect 37996 39778 38052 39788
rect 38332 39844 38388 40350
rect 38668 40178 38724 41020
rect 38780 40404 38836 41134
rect 38780 40338 38836 40348
rect 38668 40126 38670 40178
rect 38722 40126 38724 40178
rect 38668 40114 38724 40126
rect 38332 39842 38612 39844
rect 38332 39790 38334 39842
rect 38386 39790 38612 39842
rect 38332 39788 38612 39790
rect 38332 39778 38388 39788
rect 38556 38834 38612 39788
rect 38556 38782 38558 38834
rect 38610 38782 38612 38834
rect 38332 38724 38388 38762
rect 38332 38658 38388 38668
rect 37884 37998 37886 38050
rect 37938 37998 37940 38050
rect 37884 37986 37940 37998
rect 38108 38050 38164 38062
rect 38108 37998 38110 38050
rect 38162 37998 38164 38050
rect 37884 37828 37940 37838
rect 37884 37734 37940 37772
rect 38108 37380 38164 37998
rect 38108 37314 38164 37324
rect 38444 37380 38500 37390
rect 38444 37286 38500 37324
rect 38332 37266 38388 37278
rect 38332 37214 38334 37266
rect 38386 37214 38388 37266
rect 37772 36540 38164 36596
rect 37996 36370 38052 36382
rect 37996 36318 37998 36370
rect 38050 36318 38052 36370
rect 37436 35812 37492 35822
rect 37436 35718 37492 35756
rect 37548 35700 37604 35710
rect 37548 35606 37604 35644
rect 37996 35364 38052 36318
rect 38108 36260 38164 36540
rect 38332 36484 38388 37214
rect 38556 36820 38612 38782
rect 38556 36764 38836 36820
rect 38332 36428 38500 36484
rect 38108 36258 38276 36260
rect 38108 36206 38110 36258
rect 38162 36206 38276 36258
rect 38108 36204 38276 36206
rect 38108 36194 38164 36204
rect 37996 35298 38052 35308
rect 38108 35812 38164 35822
rect 37380 35196 37492 35252
rect 37324 35186 37380 35196
rect 37324 34916 37380 34926
rect 37324 34822 37380 34860
rect 37212 34750 37214 34802
rect 37266 34750 37268 34802
rect 37212 34738 37268 34750
rect 37436 33570 37492 35196
rect 38108 35028 38164 35756
rect 37884 35026 38164 35028
rect 37884 34974 38110 35026
rect 38162 34974 38164 35026
rect 37884 34972 38164 34974
rect 37884 34130 37940 34972
rect 38108 34962 38164 34972
rect 37884 34078 37886 34130
rect 37938 34078 37940 34130
rect 37884 34066 37940 34078
rect 38220 34914 38276 36204
rect 38332 36258 38388 36270
rect 38332 36206 38334 36258
rect 38386 36206 38388 36258
rect 38332 35698 38388 36206
rect 38332 35646 38334 35698
rect 38386 35646 38388 35698
rect 38332 35634 38388 35646
rect 38220 34862 38222 34914
rect 38274 34862 38276 34914
rect 38220 33908 38276 34862
rect 38220 33842 38276 33852
rect 37436 33518 37438 33570
rect 37490 33518 37492 33570
rect 37436 33506 37492 33518
rect 38220 33460 38276 33470
rect 38108 33404 38220 33460
rect 37996 33122 38052 33134
rect 37996 33070 37998 33122
rect 38050 33070 38052 33122
rect 37548 33012 37604 33022
rect 36652 32786 36708 32798
rect 36652 32734 36654 32786
rect 36706 32734 36708 32786
rect 36652 32676 36708 32734
rect 37212 32788 37268 32798
rect 37212 32694 37268 32732
rect 36652 32610 36708 32620
rect 37324 32676 37380 32686
rect 37212 32564 37268 32574
rect 37100 31892 37156 31902
rect 37212 31892 37268 32508
rect 37100 31890 37268 31892
rect 37100 31838 37102 31890
rect 37154 31838 37268 31890
rect 37100 31836 37268 31838
rect 37100 31826 37156 31836
rect 36540 31154 36596 31164
rect 33516 30942 33518 30994
rect 33570 30942 33572 30994
rect 33516 30930 33572 30942
rect 33628 31108 33684 31118
rect 33628 30996 33684 31052
rect 33964 31108 34020 31118
rect 33852 30996 33908 31006
rect 33628 30994 33908 30996
rect 33628 30942 33854 30994
rect 33906 30942 33908 30994
rect 33628 30940 33908 30942
rect 33852 30930 33908 30940
rect 33964 30212 34020 31052
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 33964 30118 34020 30156
rect 33180 29374 33182 29426
rect 33234 29374 33236 29426
rect 33180 29362 33236 29374
rect 33292 30100 33348 30110
rect 33292 28868 33348 30044
rect 33404 29986 33460 29998
rect 33628 29988 33684 29998
rect 33404 29934 33406 29986
rect 33458 29934 33460 29986
rect 33404 29652 33460 29934
rect 33404 29586 33460 29596
rect 33516 29986 33684 29988
rect 33516 29934 33630 29986
rect 33682 29934 33684 29986
rect 33516 29932 33684 29934
rect 33292 28802 33348 28812
rect 33068 28702 33070 28754
rect 33122 28702 33124 28754
rect 33068 28690 33124 28702
rect 33180 28756 33236 28766
rect 33180 28530 33236 28700
rect 33516 28642 33572 29932
rect 33628 29922 33684 29932
rect 37324 29986 37380 32620
rect 37548 32564 37604 32956
rect 37772 32676 37828 32686
rect 37996 32676 38052 33070
rect 37828 32620 38052 32676
rect 38108 32788 38164 33404
rect 38220 33394 38276 33404
rect 38108 32674 38164 32732
rect 38108 32622 38110 32674
rect 38162 32622 38164 32674
rect 37772 32582 37828 32620
rect 38108 32610 38164 32622
rect 38444 32674 38500 36428
rect 38780 35700 38836 36764
rect 38780 35606 38836 35644
rect 38668 35586 38724 35598
rect 38668 35534 38670 35586
rect 38722 35534 38724 35586
rect 38668 35364 38724 35534
rect 38668 35298 38724 35308
rect 38556 34804 38612 34814
rect 38556 34710 38612 34748
rect 38892 34354 38948 42476
rect 39004 42466 39060 42476
rect 39116 39620 39172 45724
rect 39228 45780 39284 45790
rect 39228 45686 39284 45724
rect 39340 45444 39396 45454
rect 39228 45388 39340 45444
rect 39228 44434 39284 45388
rect 39340 45378 39396 45388
rect 39228 44382 39230 44434
rect 39282 44382 39284 44434
rect 39228 44370 39284 44382
rect 39340 44434 39396 44446
rect 39340 44382 39342 44434
rect 39394 44382 39396 44434
rect 39340 43316 39396 44382
rect 39676 44322 39732 47404
rect 40236 47394 40292 47406
rect 40124 46900 40180 46910
rect 40124 46806 40180 46844
rect 40348 46898 40404 47964
rect 40348 46846 40350 46898
rect 40402 46846 40404 46898
rect 40348 46834 40404 46846
rect 39900 46786 39956 46798
rect 39900 46734 39902 46786
rect 39954 46734 39956 46786
rect 39900 46676 39956 46734
rect 40236 46676 40292 46686
rect 39900 46610 39956 46620
rect 40124 46674 40292 46676
rect 40124 46622 40238 46674
rect 40290 46622 40292 46674
rect 40124 46620 40292 46622
rect 40012 45780 40068 45790
rect 39676 44270 39678 44322
rect 39730 44270 39732 44322
rect 39676 43540 39732 44270
rect 39676 43474 39732 43484
rect 39788 45668 39844 45678
rect 39340 43250 39396 43260
rect 39788 41972 39844 45612
rect 40012 45218 40068 45724
rect 40012 45166 40014 45218
rect 40066 45166 40068 45218
rect 40012 45154 40068 45166
rect 40124 44772 40180 46620
rect 40236 46610 40292 46620
rect 40572 45332 40628 48748
rect 40908 48354 40964 48972
rect 41020 49026 41076 49038
rect 41020 48974 41022 49026
rect 41074 48974 41076 49026
rect 41020 48466 41076 48974
rect 41020 48414 41022 48466
rect 41074 48414 41076 48466
rect 41020 48402 41076 48414
rect 40908 48302 40910 48354
rect 40962 48302 40964 48354
rect 40796 48020 40852 48030
rect 40796 47458 40852 47964
rect 40796 47406 40798 47458
rect 40850 47406 40852 47458
rect 40796 47124 40852 47406
rect 40908 47346 40964 48302
rect 41244 48244 41300 48254
rect 41804 48244 41860 52780
rect 42476 52388 42532 53564
rect 43148 53620 43204 53630
rect 43148 53526 43204 53564
rect 43260 53618 43316 53676
rect 43260 53566 43262 53618
rect 43314 53566 43316 53618
rect 43260 53554 43316 53566
rect 42476 52322 42532 52332
rect 43932 52388 43988 54574
rect 45052 54516 45108 55244
rect 45276 55298 45332 55310
rect 45276 55246 45278 55298
rect 45330 55246 45332 55298
rect 45164 54516 45220 54526
rect 45052 54514 45220 54516
rect 45052 54462 45166 54514
rect 45218 54462 45220 54514
rect 45052 54460 45220 54462
rect 45164 54450 45220 54460
rect 44492 54404 44548 54414
rect 44492 54310 44548 54348
rect 44940 54402 44996 54414
rect 44940 54350 44942 54402
rect 44994 54350 44996 54402
rect 44940 54292 44996 54350
rect 45276 54292 45332 55246
rect 45836 55188 45892 55198
rect 46172 55188 46228 55198
rect 45836 55186 46228 55188
rect 45836 55134 45838 55186
rect 45890 55134 46174 55186
rect 46226 55134 46228 55186
rect 45836 55132 46228 55134
rect 45836 55122 45892 55132
rect 46172 55122 46228 55132
rect 46508 55186 46564 56028
rect 47404 56084 47460 56094
rect 47404 55990 47460 56028
rect 52444 55970 52500 59200
rect 54460 56642 54516 59200
rect 54460 56590 54462 56642
rect 54514 56590 54516 56642
rect 54460 56578 54516 56590
rect 55020 56642 55076 56654
rect 55020 56590 55022 56642
rect 55074 56590 55076 56642
rect 55020 56306 55076 56590
rect 55020 56254 55022 56306
rect 55074 56254 55076 56306
rect 55020 56242 55076 56254
rect 55132 56308 55188 59200
rect 55468 56308 55524 56318
rect 55132 56306 55524 56308
rect 55132 56254 55470 56306
rect 55522 56254 55524 56306
rect 55132 56252 55524 56254
rect 55468 56242 55524 56252
rect 52444 55918 52446 55970
rect 52498 55918 52500 55970
rect 52444 55906 52500 55918
rect 53004 56084 53060 56094
rect 46508 55134 46510 55186
rect 46562 55134 46564 55186
rect 46508 55122 46564 55134
rect 47964 55410 48020 55422
rect 47964 55358 47966 55410
rect 48018 55358 48020 55410
rect 47404 55076 47460 55086
rect 47404 55074 47572 55076
rect 47404 55022 47406 55074
rect 47458 55022 47572 55074
rect 47404 55020 47572 55022
rect 47404 55010 47460 55020
rect 45500 54740 45556 54750
rect 45500 54646 45556 54684
rect 46396 54628 46452 54638
rect 46396 54514 46452 54572
rect 46956 54628 47012 54638
rect 46956 54534 47012 54572
rect 46396 54462 46398 54514
rect 46450 54462 46452 54514
rect 46396 54450 46452 54462
rect 46844 54514 46900 54526
rect 46844 54462 46846 54514
rect 46898 54462 46900 54514
rect 44996 54236 45332 54292
rect 44940 54226 44996 54236
rect 46844 53956 46900 54462
rect 46844 53890 46900 53900
rect 47068 54514 47124 54526
rect 47068 54462 47070 54514
rect 47122 54462 47124 54514
rect 46508 53844 46564 53854
rect 45836 53732 45892 53742
rect 45724 52834 45780 52846
rect 45724 52782 45726 52834
rect 45778 52782 45780 52834
rect 45724 52724 45780 52782
rect 43932 52322 43988 52332
rect 45276 52668 45780 52724
rect 43260 52276 43316 52286
rect 43484 52276 43540 52286
rect 43260 52182 43316 52220
rect 43372 52220 43484 52276
rect 43260 52052 43316 52062
rect 42700 51940 42756 51950
rect 42476 51716 42532 51726
rect 42476 50596 42532 51660
rect 42700 51490 42756 51884
rect 42700 51438 42702 51490
rect 42754 51438 42756 51490
rect 42700 51044 42756 51438
rect 43036 51490 43092 51502
rect 43036 51438 43038 51490
rect 43090 51438 43092 51490
rect 43036 51156 43092 51438
rect 43036 51090 43092 51100
rect 43260 51156 43316 51996
rect 43372 51492 43428 52220
rect 43484 52210 43540 52220
rect 44044 52276 44100 52286
rect 44044 52182 44100 52220
rect 45164 52276 45220 52286
rect 43596 52164 43652 52174
rect 43596 52070 43652 52108
rect 43820 52162 43876 52174
rect 43820 52110 43822 52162
rect 43874 52110 43876 52162
rect 43484 52052 43540 52062
rect 43484 51958 43540 51996
rect 43372 51436 43652 51492
rect 43484 51268 43540 51278
rect 43372 51266 43540 51268
rect 43372 51214 43486 51266
rect 43538 51214 43540 51266
rect 43372 51212 43540 51214
rect 43372 51156 43428 51212
rect 43484 51202 43540 51212
rect 43260 51100 43428 51156
rect 42700 50978 42756 50988
rect 42252 50594 42532 50596
rect 42252 50542 42478 50594
rect 42530 50542 42532 50594
rect 42252 50540 42532 50542
rect 42140 50482 42196 50494
rect 42140 50430 42142 50482
rect 42194 50430 42196 50482
rect 42140 50260 42196 50430
rect 42140 50194 42196 50204
rect 42140 49812 42196 49822
rect 42252 49812 42308 50540
rect 42476 50530 42532 50540
rect 43260 50596 43316 51100
rect 43484 51044 43540 51054
rect 42812 50372 42868 50382
rect 42812 50278 42868 50316
rect 42140 49810 42308 49812
rect 42140 49758 42142 49810
rect 42194 49758 42308 49810
rect 42140 49756 42308 49758
rect 42140 49746 42196 49756
rect 43260 48468 43316 50540
rect 43372 50594 43428 50606
rect 43372 50542 43374 50594
rect 43426 50542 43428 50594
rect 43372 50260 43428 50542
rect 43372 49924 43428 50204
rect 43372 49858 43428 49868
rect 43484 49922 43540 50988
rect 43484 49870 43486 49922
rect 43538 49870 43540 49922
rect 43484 49858 43540 49870
rect 43596 50372 43652 51436
rect 43708 51156 43764 51166
rect 43820 51156 43876 52110
rect 44828 52164 44884 52174
rect 44828 52070 44884 52108
rect 45052 52052 45108 52062
rect 44940 52050 45108 52052
rect 44940 51998 45054 52050
rect 45106 51998 45108 52050
rect 44940 51996 45108 51998
rect 45164 52052 45220 52220
rect 45276 52274 45332 52668
rect 45276 52222 45278 52274
rect 45330 52222 45332 52274
rect 45276 52210 45332 52222
rect 45612 52500 45668 52510
rect 45388 52052 45444 52062
rect 45164 52050 45444 52052
rect 45164 51998 45390 52050
rect 45442 51998 45444 52050
rect 45164 51996 45444 51998
rect 44940 51716 44996 51996
rect 45052 51986 45108 51996
rect 45388 51986 45444 51996
rect 44044 51660 44996 51716
rect 44044 51602 44100 51660
rect 44044 51550 44046 51602
rect 44098 51550 44100 51602
rect 44044 51538 44100 51550
rect 43764 51100 43876 51156
rect 43708 51062 43764 51100
rect 43596 48916 43652 50316
rect 43708 50706 43764 50718
rect 43708 50654 43710 50706
rect 43762 50654 43764 50706
rect 43708 49138 43764 50654
rect 43708 49086 43710 49138
rect 43762 49086 43764 49138
rect 43708 49074 43764 49086
rect 43820 49028 43876 51100
rect 45612 50596 45668 52444
rect 45724 52162 45780 52668
rect 45836 52386 45892 53676
rect 46508 53058 46564 53788
rect 47068 53844 47124 54462
rect 47068 53778 47124 53788
rect 47404 54402 47460 54414
rect 47404 54350 47406 54402
rect 47458 54350 47460 54402
rect 47180 53732 47236 53742
rect 47180 53638 47236 53676
rect 46508 53006 46510 53058
rect 46562 53006 46564 53058
rect 46508 52994 46564 53006
rect 45836 52334 45838 52386
rect 45890 52334 45892 52386
rect 45836 52322 45892 52334
rect 45948 52946 46004 52958
rect 45948 52894 45950 52946
rect 46002 52894 46004 52946
rect 45724 52110 45726 52162
rect 45778 52110 45780 52162
rect 45724 52098 45780 52110
rect 45836 51940 45892 51950
rect 45948 51940 46004 52894
rect 45836 51938 46004 51940
rect 45836 51886 45838 51938
rect 45890 51886 46004 51938
rect 45836 51884 46004 51886
rect 46172 52388 46228 52398
rect 45836 51268 45892 51884
rect 46172 51492 46228 52332
rect 47404 52276 47460 54350
rect 47516 53956 47572 55020
rect 47628 54516 47684 54526
rect 47964 54516 48020 55358
rect 51212 55298 51268 55310
rect 51212 55246 51214 55298
rect 51266 55246 51268 55298
rect 48188 55186 48244 55198
rect 48188 55134 48190 55186
rect 48242 55134 48244 55186
rect 48188 55076 48244 55134
rect 49868 55188 49924 55198
rect 49868 55186 50036 55188
rect 49868 55134 49870 55186
rect 49922 55134 50036 55186
rect 49868 55132 50036 55134
rect 49868 55122 49924 55132
rect 48188 55010 48244 55020
rect 48748 55076 48804 55086
rect 47684 54460 48020 54516
rect 47628 54422 47684 54460
rect 47516 53890 47572 53900
rect 47852 54292 47908 54302
rect 47740 53844 47796 53854
rect 47852 53844 47908 54236
rect 47796 53788 47908 53844
rect 47740 53730 47796 53788
rect 47740 53678 47742 53730
rect 47794 53678 47796 53730
rect 47740 53666 47796 53678
rect 47964 53730 48020 54460
rect 48300 54516 48356 54526
rect 48300 54422 48356 54460
rect 48748 54514 48804 55020
rect 49980 54738 50036 55132
rect 50764 55076 50820 55086
rect 51212 55076 51268 55246
rect 50764 55074 51268 55076
rect 50764 55022 50766 55074
rect 50818 55022 51268 55074
rect 50764 55020 51268 55022
rect 50764 55010 50820 55020
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 49980 54686 49982 54738
rect 50034 54686 50036 54738
rect 49980 54674 50036 54686
rect 50764 54740 50820 54750
rect 49084 54628 49140 54638
rect 49084 54534 49140 54572
rect 50764 54626 50820 54684
rect 50764 54574 50766 54626
rect 50818 54574 50820 54626
rect 50764 54562 50820 54574
rect 48748 54462 48750 54514
rect 48802 54462 48804 54514
rect 48748 54450 48804 54462
rect 48972 54516 49028 54526
rect 48972 54422 49028 54460
rect 49532 54516 49588 54526
rect 49532 54422 49588 54460
rect 50204 54514 50260 54526
rect 50204 54462 50206 54514
rect 50258 54462 50260 54514
rect 49196 54404 49252 54414
rect 49252 54348 49364 54404
rect 49196 54338 49252 54348
rect 47964 53678 47966 53730
rect 48018 53678 48020 53730
rect 47964 53666 48020 53678
rect 48076 53956 48132 53966
rect 47628 53620 47684 53630
rect 47628 53526 47684 53564
rect 47404 52210 47460 52220
rect 45836 51202 45892 51212
rect 45948 51490 46228 51492
rect 45948 51438 46174 51490
rect 46226 51438 46228 51490
rect 45948 51436 46228 51438
rect 45948 50708 46004 51436
rect 46172 51426 46228 51436
rect 46732 51938 46788 51950
rect 46732 51886 46734 51938
rect 46786 51886 46788 51938
rect 46508 51268 46564 51278
rect 46732 51268 46788 51886
rect 47180 51940 47236 51950
rect 47628 51940 47684 51950
rect 47180 51938 47684 51940
rect 47180 51886 47182 51938
rect 47234 51886 47630 51938
rect 47682 51886 47684 51938
rect 47180 51884 47684 51886
rect 47180 51874 47236 51884
rect 47068 51604 47124 51614
rect 47124 51548 47236 51604
rect 47068 51538 47124 51548
rect 46956 51268 47012 51278
rect 46732 51212 46956 51268
rect 46508 51174 46564 51212
rect 46956 51174 47012 51212
rect 45612 50502 45668 50540
rect 45724 50652 46004 50708
rect 44268 50484 44324 50494
rect 44268 50390 44324 50428
rect 44380 50036 44436 50046
rect 44380 49924 44436 49980
rect 45276 49924 45332 49934
rect 44380 49922 44884 49924
rect 44380 49870 44382 49922
rect 44434 49870 44884 49922
rect 44380 49868 44884 49870
rect 44380 49858 44436 49868
rect 43820 48934 43876 48972
rect 44268 49252 44324 49262
rect 43596 48822 43652 48860
rect 44156 48914 44212 48926
rect 44156 48862 44158 48914
rect 44210 48862 44212 48914
rect 43484 48468 43540 48478
rect 43260 48466 43764 48468
rect 43260 48414 43486 48466
rect 43538 48414 43764 48466
rect 43260 48412 43764 48414
rect 43484 48402 43540 48412
rect 41244 48242 41636 48244
rect 41244 48190 41246 48242
rect 41298 48190 41636 48242
rect 41244 48188 41636 48190
rect 41804 48188 42084 48244
rect 41244 48178 41300 48188
rect 40908 47294 40910 47346
rect 40962 47294 40964 47346
rect 40908 47282 40964 47294
rect 41244 47570 41300 47582
rect 41244 47518 41246 47570
rect 41298 47518 41300 47570
rect 40796 47068 41076 47124
rect 41020 46786 41076 47068
rect 41020 46734 41022 46786
rect 41074 46734 41076 46786
rect 41020 46722 41076 46734
rect 40908 46676 40964 46686
rect 40908 46582 40964 46620
rect 41244 46676 41300 47518
rect 41244 46610 41300 46620
rect 41580 47348 41636 48188
rect 41692 48132 41748 48142
rect 41692 48130 41972 48132
rect 41692 48078 41694 48130
rect 41746 48078 41972 48130
rect 41692 48076 41972 48078
rect 41692 48066 41748 48076
rect 41916 47458 41972 48076
rect 41916 47406 41918 47458
rect 41970 47406 41972 47458
rect 41692 47348 41748 47358
rect 41580 47346 41860 47348
rect 41580 47294 41694 47346
rect 41746 47294 41860 47346
rect 41580 47292 41860 47294
rect 41580 46900 41636 47292
rect 41692 47282 41748 47292
rect 41468 46562 41524 46574
rect 41468 46510 41470 46562
rect 41522 46510 41524 46562
rect 41244 46116 41300 46126
rect 41244 46022 41300 46060
rect 40124 44706 40180 44716
rect 40236 45276 40628 45332
rect 41356 45666 41412 45678
rect 41356 45614 41358 45666
rect 41410 45614 41412 45666
rect 40236 44660 40292 45276
rect 40348 45108 40404 45118
rect 40348 45106 40964 45108
rect 40348 45054 40350 45106
rect 40402 45054 40964 45106
rect 40348 45052 40964 45054
rect 40348 45042 40404 45052
rect 40908 44996 40964 45052
rect 41356 45106 41412 45614
rect 41356 45054 41358 45106
rect 41410 45054 41412 45106
rect 41356 45042 41412 45054
rect 40908 44940 41300 44996
rect 40348 44884 40404 44894
rect 40348 44882 40852 44884
rect 40348 44830 40350 44882
rect 40402 44830 40852 44882
rect 40348 44828 40852 44830
rect 40348 44818 40404 44828
rect 40236 44604 40516 44660
rect 40348 43540 40404 43550
rect 39228 41970 39844 41972
rect 39228 41918 39790 41970
rect 39842 41918 39844 41970
rect 39228 41916 39844 41918
rect 39228 41186 39284 41916
rect 39788 41906 39844 41916
rect 40236 41972 40292 41982
rect 40236 41858 40292 41916
rect 40236 41806 40238 41858
rect 40290 41806 40292 41858
rect 40236 41794 40292 41806
rect 39228 41134 39230 41186
rect 39282 41134 39284 41186
rect 39228 41122 39284 41134
rect 39676 41188 39732 41198
rect 39676 41094 39732 41132
rect 39564 39620 39620 39630
rect 39116 39618 39620 39620
rect 39116 39566 39566 39618
rect 39618 39566 39620 39618
rect 39116 39564 39620 39566
rect 39564 39554 39620 39564
rect 39900 39396 39956 39406
rect 39900 39302 39956 39340
rect 39228 38724 39284 38762
rect 39228 38658 39284 38668
rect 39004 37828 39060 37838
rect 39004 37266 39060 37772
rect 39004 37214 39006 37266
rect 39058 37214 39060 37266
rect 39004 37202 39060 37214
rect 39116 37492 39172 37502
rect 39116 36370 39172 37436
rect 39788 37492 39844 37502
rect 39340 37380 39396 37390
rect 39340 37286 39396 37324
rect 39788 37266 39844 37436
rect 40348 37490 40404 43484
rect 40460 41300 40516 44604
rect 40796 44322 40852 44828
rect 40796 44270 40798 44322
rect 40850 44270 40852 44322
rect 40796 44258 40852 44270
rect 41020 44772 41076 44782
rect 41020 44322 41076 44716
rect 41020 44270 41022 44322
rect 41074 44270 41076 44322
rect 41020 44258 41076 44270
rect 41244 44322 41300 44940
rect 41356 44548 41412 44558
rect 41468 44548 41524 46510
rect 41580 45890 41636 46844
rect 41804 46674 41860 47292
rect 41916 47012 41972 47406
rect 41916 46946 41972 46956
rect 42028 46788 42084 48188
rect 43708 47458 43764 48412
rect 43708 47406 43710 47458
rect 43762 47406 43764 47458
rect 43708 47394 43764 47406
rect 43820 48242 43876 48254
rect 43820 48190 43822 48242
rect 43874 48190 43876 48242
rect 43820 48132 43876 48190
rect 44156 48132 44212 48862
rect 43820 48130 44212 48132
rect 43820 48078 44158 48130
rect 44210 48078 44212 48130
rect 43820 48076 44212 48078
rect 41804 46622 41806 46674
rect 41858 46622 41860 46674
rect 41804 46610 41860 46622
rect 41916 46732 42084 46788
rect 41580 45838 41582 45890
rect 41634 45838 41636 45890
rect 41580 45826 41636 45838
rect 41916 45780 41972 46732
rect 42252 46676 42308 46686
rect 41916 45714 41972 45724
rect 42140 46116 42196 46126
rect 42028 45218 42084 45230
rect 42028 45166 42030 45218
rect 42082 45166 42084 45218
rect 41804 44994 41860 45006
rect 41804 44942 41806 44994
rect 41858 44942 41860 44994
rect 41468 44492 41636 44548
rect 41356 44434 41412 44492
rect 41356 44382 41358 44434
rect 41410 44382 41412 44434
rect 41356 44370 41412 44382
rect 41244 44270 41246 44322
rect 41298 44270 41300 44322
rect 41244 43764 41300 44270
rect 41468 44322 41524 44334
rect 41468 44270 41470 44322
rect 41522 44270 41524 44322
rect 41468 44100 41524 44270
rect 41468 44034 41524 44044
rect 41244 43762 41412 43764
rect 41244 43710 41246 43762
rect 41298 43710 41412 43762
rect 41244 43708 41412 43710
rect 41244 43698 41300 43708
rect 40908 43540 40964 43550
rect 40908 43446 40964 43484
rect 41356 42754 41412 43708
rect 41356 42702 41358 42754
rect 41410 42702 41412 42754
rect 41356 42194 41412 42702
rect 41356 42142 41358 42194
rect 41410 42142 41412 42194
rect 41356 42130 41412 42142
rect 41580 41300 41636 44492
rect 41804 43540 41860 44942
rect 41804 43474 41860 43484
rect 42028 44100 42084 45166
rect 42140 45106 42196 46060
rect 42140 45054 42142 45106
rect 42194 45054 42196 45106
rect 42140 45042 42196 45054
rect 41916 42754 41972 42766
rect 41916 42702 41918 42754
rect 41970 42702 41972 42754
rect 41916 42644 41972 42702
rect 41916 42578 41972 42588
rect 42028 41972 42084 44044
rect 42252 42754 42308 46620
rect 42476 46674 42532 46686
rect 42476 46622 42478 46674
rect 42530 46622 42532 46674
rect 42476 45444 42532 46622
rect 42924 46676 42980 46686
rect 42924 46582 42980 46620
rect 42476 45378 42532 45388
rect 43372 45220 43428 45230
rect 43372 44546 43428 45164
rect 43372 44494 43374 44546
rect 43426 44494 43428 44546
rect 43372 44482 43428 44494
rect 43484 44884 43540 44894
rect 43484 44546 43540 44828
rect 43484 44494 43486 44546
rect 43538 44494 43540 44546
rect 43484 44482 43540 44494
rect 42700 44324 42756 44334
rect 43148 44324 43204 44334
rect 42756 44322 43204 44324
rect 42756 44270 43150 44322
rect 43202 44270 43204 44322
rect 42756 44268 43204 44270
rect 42700 44230 42756 44268
rect 43148 44258 43204 44268
rect 43484 44100 43540 44110
rect 43484 44006 43540 44044
rect 42588 43540 42644 43550
rect 42588 43446 42644 43484
rect 42924 43540 42980 43550
rect 43708 43540 43764 43550
rect 42924 42868 42980 43484
rect 43596 43538 43764 43540
rect 43596 43486 43710 43538
rect 43762 43486 43764 43538
rect 43596 43484 43764 43486
rect 42252 42702 42254 42754
rect 42306 42702 42308 42754
rect 42028 41906 42084 41916
rect 42140 41970 42196 41982
rect 42140 41918 42142 41970
rect 42194 41918 42196 41970
rect 40460 41298 40964 41300
rect 40460 41246 40462 41298
rect 40514 41246 40964 41298
rect 40460 41244 40964 41246
rect 40460 41234 40516 41244
rect 40348 37438 40350 37490
rect 40402 37438 40404 37490
rect 40348 37426 40404 37438
rect 40908 41186 40964 41244
rect 40908 41134 40910 41186
rect 40962 41134 40964 41186
rect 39788 37214 39790 37266
rect 39842 37214 39844 37266
rect 39788 37202 39844 37214
rect 40012 37042 40068 37054
rect 40012 36990 40014 37042
rect 40066 36990 40068 37042
rect 39116 36318 39118 36370
rect 39170 36318 39172 36370
rect 39116 34914 39172 36318
rect 39116 34862 39118 34914
rect 39170 34862 39172 34914
rect 39116 34850 39172 34862
rect 39340 36484 39396 36494
rect 40012 36484 40068 36990
rect 39340 36482 40068 36484
rect 39340 36430 39342 36482
rect 39394 36430 40068 36482
rect 39340 36428 40068 36430
rect 38892 34302 38894 34354
rect 38946 34302 38948 34354
rect 38892 34290 38948 34302
rect 39228 34242 39284 34254
rect 39228 34190 39230 34242
rect 39282 34190 39284 34242
rect 38668 34130 38724 34142
rect 38668 34078 38670 34130
rect 38722 34078 38724 34130
rect 38668 33460 38724 34078
rect 39228 33572 39284 34190
rect 39228 33506 39284 33516
rect 38668 33394 38724 33404
rect 38444 32622 38446 32674
rect 38498 32622 38500 32674
rect 37548 32470 37604 32508
rect 38444 31948 38500 32622
rect 38444 31892 38724 31948
rect 38332 31220 38388 31230
rect 37324 29934 37326 29986
rect 37378 29934 37380 29986
rect 36316 29652 36372 29662
rect 36316 29558 36372 29596
rect 37324 29652 37380 29934
rect 37660 29988 37716 29998
rect 38332 29988 38388 31164
rect 38556 31218 38612 31892
rect 38668 31780 38724 31892
rect 38668 31686 38724 31724
rect 39004 31890 39060 31902
rect 39004 31838 39006 31890
rect 39058 31838 39060 31890
rect 38556 31166 38558 31218
rect 38610 31166 38612 31218
rect 38556 31154 38612 31166
rect 38780 31220 38836 31230
rect 38780 31126 38836 31164
rect 39004 31220 39060 31838
rect 39340 31890 39396 36428
rect 39564 36260 39620 36270
rect 39564 36166 39620 36204
rect 40908 36260 40964 41134
rect 41132 41244 41636 41300
rect 41132 41074 41188 41244
rect 41132 41022 41134 41074
rect 41186 41022 41188 41074
rect 41132 41010 41188 41022
rect 41580 39172 41636 41244
rect 41916 41858 41972 41870
rect 41916 41806 41918 41858
rect 41970 41806 41972 41858
rect 41692 41188 41748 41198
rect 41692 40626 41748 41132
rect 41692 40574 41694 40626
rect 41746 40574 41748 40626
rect 41692 40562 41748 40574
rect 41804 40628 41860 40638
rect 41804 40534 41860 40572
rect 41916 40626 41972 41806
rect 42028 41412 42084 41422
rect 42028 41318 42084 41356
rect 41916 40574 41918 40626
rect 41970 40574 41972 40626
rect 41916 39956 41972 40574
rect 42140 40626 42196 41918
rect 42140 40574 42142 40626
rect 42194 40574 42196 40626
rect 42140 40562 42196 40574
rect 41916 39900 42196 39956
rect 42140 39620 42196 39900
rect 42252 39844 42308 42702
rect 42812 42866 42980 42868
rect 42812 42814 42926 42866
rect 42978 42814 42980 42866
rect 42812 42812 42980 42814
rect 42588 42644 42644 42654
rect 42364 42588 42588 42644
rect 42364 42194 42420 42588
rect 42588 42550 42644 42588
rect 42364 42142 42366 42194
rect 42418 42142 42420 42194
rect 42364 42130 42420 42142
rect 42476 41972 42532 41982
rect 42476 41300 42532 41916
rect 42588 41300 42644 41310
rect 42476 41298 42644 41300
rect 42476 41246 42590 41298
rect 42642 41246 42644 41298
rect 42476 41244 42644 41246
rect 42588 41234 42644 41244
rect 42364 39844 42420 39854
rect 42252 39842 42420 39844
rect 42252 39790 42366 39842
rect 42418 39790 42420 39842
rect 42252 39788 42420 39790
rect 42364 39778 42420 39788
rect 42140 39618 42308 39620
rect 42140 39566 42142 39618
rect 42194 39566 42308 39618
rect 42140 39564 42308 39566
rect 42140 39554 42196 39564
rect 41580 39106 41636 39116
rect 41804 39396 41860 39406
rect 42252 39396 42308 39564
rect 42700 39396 42756 39406
rect 42252 39340 42532 39396
rect 41804 38946 41860 39340
rect 41804 38894 41806 38946
rect 41858 38894 41860 38946
rect 41580 38836 41636 38846
rect 41580 38276 41636 38780
rect 41580 38210 41636 38220
rect 41356 37940 41412 37950
rect 41020 37716 41076 37726
rect 41020 37266 41076 37660
rect 41356 37490 41412 37884
rect 41804 37492 41860 38894
rect 42364 39172 42420 39182
rect 42140 38836 42196 38846
rect 42140 38742 42196 38780
rect 42252 37940 42308 37950
rect 42252 37846 42308 37884
rect 41356 37438 41358 37490
rect 41410 37438 41412 37490
rect 41356 37426 41412 37438
rect 41580 37436 41860 37492
rect 41020 37214 41022 37266
rect 41074 37214 41076 37266
rect 41020 37044 41076 37214
rect 41020 36978 41076 36988
rect 41356 37268 41412 37278
rect 41580 37268 41636 37436
rect 41356 37266 41636 37268
rect 41356 37214 41358 37266
rect 41410 37214 41636 37266
rect 41356 37212 41636 37214
rect 41692 37268 41748 37278
rect 42140 37268 42196 37278
rect 41692 37266 42196 37268
rect 41692 37214 41694 37266
rect 41746 37214 42142 37266
rect 42194 37214 42196 37266
rect 41692 37212 42196 37214
rect 40908 36194 40964 36204
rect 41244 36596 41300 36606
rect 39452 35810 39508 35822
rect 39452 35758 39454 35810
rect 39506 35758 39508 35810
rect 39452 35700 39508 35758
rect 41244 35810 41300 36540
rect 41244 35758 41246 35810
rect 41298 35758 41300 35810
rect 41244 35746 41300 35758
rect 41356 35810 41412 37212
rect 41692 37202 41748 37212
rect 42140 37202 42196 37212
rect 42364 37266 42420 39116
rect 42476 38834 42532 39340
rect 42700 39302 42756 39340
rect 42588 39058 42644 39070
rect 42588 39006 42590 39058
rect 42642 39006 42644 39058
rect 42588 38948 42644 39006
rect 42588 38882 42644 38892
rect 42476 38782 42478 38834
rect 42530 38782 42532 38834
rect 42476 38050 42532 38782
rect 42476 37998 42478 38050
rect 42530 37998 42532 38050
rect 42476 37986 42532 37998
rect 42812 38052 42868 42812
rect 42924 42802 42980 42812
rect 43484 43428 43540 43438
rect 42924 42644 42980 42654
rect 42924 41186 42980 42588
rect 43484 41300 43540 43372
rect 43596 42644 43652 43484
rect 43708 43474 43764 43484
rect 43596 42578 43652 42588
rect 43484 41244 43652 41300
rect 42924 41134 42926 41186
rect 42978 41134 42980 41186
rect 42924 41122 42980 41134
rect 43484 41076 43540 41086
rect 43148 41074 43540 41076
rect 43148 41022 43486 41074
rect 43538 41022 43540 41074
rect 43148 41020 43540 41022
rect 43036 39172 43092 39182
rect 43036 38946 43092 39116
rect 43036 38894 43038 38946
rect 43090 38894 43092 38946
rect 43036 38882 43092 38894
rect 43148 38388 43204 41020
rect 43484 41010 43540 41020
rect 43596 40852 43652 41244
rect 43484 40796 43652 40852
rect 43260 38836 43316 38846
rect 43260 38742 43316 38780
rect 43036 38332 43204 38388
rect 43036 38164 43092 38332
rect 43036 38108 43204 38164
rect 42812 37986 42868 37996
rect 42364 37214 42366 37266
rect 42418 37214 42420 37266
rect 42028 37044 42084 37054
rect 42028 36950 42084 36988
rect 41804 36596 41860 36606
rect 41804 36502 41860 36540
rect 41580 36482 41636 36494
rect 41580 36430 41582 36482
rect 41634 36430 41636 36482
rect 41580 35922 41636 36430
rect 42252 36484 42308 36494
rect 42364 36484 42420 37214
rect 42252 36482 42420 36484
rect 42252 36430 42254 36482
rect 42306 36430 42420 36482
rect 42252 36428 42420 36430
rect 42252 36418 42308 36428
rect 42588 36370 42644 36382
rect 42588 36318 42590 36370
rect 42642 36318 42644 36370
rect 41580 35870 41582 35922
rect 41634 35870 41636 35922
rect 41580 35858 41636 35870
rect 42364 36260 42420 36270
rect 42364 35922 42420 36204
rect 42364 35870 42366 35922
rect 42418 35870 42420 35922
rect 42364 35858 42420 35870
rect 41356 35758 41358 35810
rect 41410 35758 41412 35810
rect 39452 35634 39508 35644
rect 41356 35588 41412 35758
rect 42588 35700 42644 36318
rect 43036 36260 43092 36270
rect 43036 35810 43092 36204
rect 43036 35758 43038 35810
rect 43090 35758 43092 35810
rect 43036 35746 43092 35758
rect 42812 35700 42868 35710
rect 42588 35698 42868 35700
rect 42588 35646 42814 35698
rect 42866 35646 42868 35698
rect 42588 35644 42868 35646
rect 42812 35634 42868 35644
rect 41244 35532 41412 35588
rect 40572 35028 40628 35038
rect 40572 34934 40628 34972
rect 39452 34690 39508 34702
rect 39452 34638 39454 34690
rect 39506 34638 39508 34690
rect 39452 34244 39508 34638
rect 40012 34244 40068 34254
rect 39452 34242 40068 34244
rect 39452 34190 40014 34242
rect 40066 34190 40068 34242
rect 39452 34188 40068 34190
rect 39452 34130 39508 34188
rect 40012 34178 40068 34188
rect 40348 34242 40404 34254
rect 40348 34190 40350 34242
rect 40402 34190 40404 34242
rect 39452 34078 39454 34130
rect 39506 34078 39508 34130
rect 39452 34066 39508 34078
rect 40348 34132 40404 34190
rect 41020 34132 41076 34142
rect 40348 34130 41076 34132
rect 40348 34078 41022 34130
rect 41074 34078 41076 34130
rect 40348 34076 41076 34078
rect 39340 31838 39342 31890
rect 39394 31838 39396 31890
rect 39340 31826 39396 31838
rect 39788 33572 39844 33582
rect 39004 31126 39060 31164
rect 39676 31220 39732 31230
rect 39788 31220 39844 33516
rect 40908 33572 40964 33582
rect 40460 33460 40516 33470
rect 40460 33346 40516 33404
rect 40460 33294 40462 33346
rect 40514 33294 40516 33346
rect 40460 33282 40516 33294
rect 40908 33346 40964 33516
rect 40908 33294 40910 33346
rect 40962 33294 40964 33346
rect 39676 31218 39844 31220
rect 39676 31166 39678 31218
rect 39730 31166 39844 31218
rect 39676 31164 39844 31166
rect 38668 30882 38724 30894
rect 38668 30830 38670 30882
rect 38722 30830 38724 30882
rect 38668 30772 38724 30830
rect 39452 30772 39508 30782
rect 38668 30770 39508 30772
rect 38668 30718 39454 30770
rect 39506 30718 39508 30770
rect 38668 30716 39508 30718
rect 39452 30706 39508 30716
rect 38892 30436 38948 30446
rect 38892 30342 38948 30380
rect 39676 30436 39732 31164
rect 40908 31106 40964 33294
rect 41020 32228 41076 34076
rect 41020 32162 41076 32172
rect 40908 31054 40910 31106
rect 40962 31054 40964 31106
rect 40908 31042 40964 31054
rect 41244 31106 41300 35532
rect 43036 35140 43092 35150
rect 43148 35140 43204 38108
rect 43372 38162 43428 38174
rect 43372 38110 43374 38162
rect 43426 38110 43428 38162
rect 43260 38052 43316 38062
rect 43260 37958 43316 37996
rect 43372 35924 43428 38110
rect 43484 38052 43540 40796
rect 43596 39060 43652 39070
rect 43596 38966 43652 39004
rect 43820 38668 43876 48076
rect 44156 48066 44212 48076
rect 44268 48466 44324 49196
rect 44268 48414 44270 48466
rect 44322 48414 44324 48466
rect 44268 47572 44324 48414
rect 44828 49138 44884 49868
rect 45276 49812 45332 49868
rect 45276 49810 45444 49812
rect 45276 49758 45278 49810
rect 45330 49758 45444 49810
rect 45276 49756 45444 49758
rect 45276 49746 45332 49756
rect 45164 49588 45220 49598
rect 45164 49586 45332 49588
rect 45164 49534 45166 49586
rect 45218 49534 45332 49586
rect 45164 49532 45332 49534
rect 45164 49522 45220 49532
rect 44828 49086 44830 49138
rect 44882 49086 44884 49138
rect 44828 48466 44884 49086
rect 44828 48414 44830 48466
rect 44882 48414 44884 48466
rect 44828 48402 44884 48414
rect 44940 48802 44996 48814
rect 44940 48750 44942 48802
rect 44994 48750 44996 48802
rect 44940 48244 44996 48750
rect 44940 48178 44996 48188
rect 45164 48354 45220 48366
rect 45164 48302 45166 48354
rect 45218 48302 45220 48354
rect 44156 47516 44324 47572
rect 44044 47124 44100 47134
rect 44044 46786 44100 47068
rect 44156 47012 44212 47516
rect 45164 47458 45220 48302
rect 45164 47406 45166 47458
rect 45218 47406 45220 47458
rect 44268 47348 44324 47358
rect 44268 47346 44772 47348
rect 44268 47294 44270 47346
rect 44322 47294 44772 47346
rect 44268 47292 44772 47294
rect 44268 47282 44324 47292
rect 44156 46946 44212 46956
rect 44044 46734 44046 46786
rect 44098 46734 44100 46786
rect 44044 46722 44100 46734
rect 44716 44324 44772 47292
rect 45164 46900 45220 47406
rect 44940 46674 44996 46686
rect 45164 46676 45220 46844
rect 44940 46622 44942 46674
rect 44994 46622 44996 46674
rect 44940 45890 44996 46622
rect 44940 45838 44942 45890
rect 44994 45838 44996 45890
rect 44940 44884 44996 45838
rect 45052 46674 45220 46676
rect 45052 46622 45166 46674
rect 45218 46622 45220 46674
rect 45052 46620 45220 46622
rect 45052 45218 45108 46620
rect 45164 46610 45220 46620
rect 45276 47012 45332 49532
rect 45388 49140 45444 49756
rect 45388 49074 45444 49084
rect 45612 49028 45668 49038
rect 45612 48914 45668 48972
rect 45612 48862 45614 48914
rect 45666 48862 45668 48914
rect 45612 48850 45668 48862
rect 45500 48802 45556 48814
rect 45500 48750 45502 48802
rect 45554 48750 45556 48802
rect 45500 48244 45556 48750
rect 45388 48242 45556 48244
rect 45388 48190 45502 48242
rect 45554 48190 45556 48242
rect 45388 48188 45556 48190
rect 45388 47458 45444 48188
rect 45500 48178 45556 48188
rect 45612 48244 45668 48254
rect 45388 47406 45390 47458
rect 45442 47406 45444 47458
rect 45388 47394 45444 47406
rect 45500 47460 45556 47470
rect 45612 47460 45668 48188
rect 45500 47458 45668 47460
rect 45500 47406 45502 47458
rect 45554 47406 45668 47458
rect 45500 47404 45668 47406
rect 45500 47394 45556 47404
rect 45276 46956 45556 47012
rect 45276 45890 45332 46956
rect 45500 46786 45556 46956
rect 45500 46734 45502 46786
rect 45554 46734 45556 46786
rect 45500 46722 45556 46734
rect 45276 45838 45278 45890
rect 45330 45838 45332 45890
rect 45276 45332 45332 45838
rect 45052 45166 45054 45218
rect 45106 45166 45108 45218
rect 45052 45154 45108 45166
rect 45164 45276 45332 45332
rect 45388 46562 45444 46574
rect 45388 46510 45390 46562
rect 45442 46510 45444 46562
rect 45164 45220 45220 45276
rect 45164 45126 45220 45164
rect 44940 44818 44996 44828
rect 45276 45106 45332 45118
rect 45276 45054 45278 45106
rect 45330 45054 45332 45106
rect 45276 44884 45332 45054
rect 45388 45108 45444 46510
rect 45500 45780 45556 45790
rect 45500 45778 45668 45780
rect 45500 45726 45502 45778
rect 45554 45726 45668 45778
rect 45500 45724 45668 45726
rect 45500 45714 45556 45724
rect 45388 45042 45444 45052
rect 45276 44818 45332 44828
rect 45052 44324 45108 44334
rect 44716 44322 45108 44324
rect 44716 44270 45054 44322
rect 45106 44270 45108 44322
rect 44716 44268 45108 44270
rect 44828 44100 44884 44110
rect 44828 44006 44884 44044
rect 44940 44098 44996 44110
rect 44940 44046 44942 44098
rect 44994 44046 44996 44098
rect 44380 43540 44436 43550
rect 44380 43446 44436 43484
rect 44940 42754 44996 44046
rect 44940 42702 44942 42754
rect 44994 42702 44996 42754
rect 44940 42690 44996 42702
rect 45052 43204 45108 44268
rect 45276 44324 45332 44334
rect 45276 43538 45332 44268
rect 45276 43486 45278 43538
rect 45330 43486 45332 43538
rect 45276 43474 45332 43486
rect 45388 44322 45444 44334
rect 45388 44270 45390 44322
rect 45442 44270 45444 44322
rect 44380 41860 44436 41870
rect 44828 41860 44884 41870
rect 44380 41858 44884 41860
rect 44380 41806 44382 41858
rect 44434 41806 44830 41858
rect 44882 41806 44884 41858
rect 44380 41804 44884 41806
rect 44380 41794 44436 41804
rect 44492 40292 44548 41804
rect 44828 41794 44884 41804
rect 44940 40292 44996 40302
rect 44492 40290 44996 40292
rect 44492 40238 44494 40290
rect 44546 40238 44942 40290
rect 44994 40238 44996 40290
rect 44492 40236 44996 40238
rect 44492 38668 44548 40236
rect 44940 40226 44996 40236
rect 45052 39956 45108 43148
rect 45276 43314 45332 43326
rect 45276 43262 45278 43314
rect 45330 43262 45332 43314
rect 45276 42756 45332 43262
rect 45388 42980 45444 44270
rect 45388 42866 45444 42924
rect 45388 42814 45390 42866
rect 45442 42814 45444 42866
rect 45388 42802 45444 42814
rect 45500 43204 45556 43214
rect 45276 42690 45332 42700
rect 45500 42754 45556 43148
rect 45500 42702 45502 42754
rect 45554 42702 45556 42754
rect 45500 42690 45556 42702
rect 45612 42084 45668 45724
rect 45724 45668 45780 50652
rect 46060 50596 46116 50606
rect 45948 50484 46004 50494
rect 45948 49810 46004 50428
rect 45948 49758 45950 49810
rect 46002 49758 46004 49810
rect 45948 49746 46004 49758
rect 46060 49588 46116 50540
rect 46172 50594 46228 50606
rect 46172 50542 46174 50594
rect 46226 50542 46228 50594
rect 46172 49924 46228 50542
rect 46284 50596 46340 50606
rect 46508 50596 46564 50606
rect 46340 50594 46564 50596
rect 46340 50542 46510 50594
rect 46562 50542 46564 50594
rect 46340 50540 46564 50542
rect 46284 50530 46340 50540
rect 46508 50530 46564 50540
rect 46732 50484 46788 50494
rect 46732 50390 46788 50428
rect 46844 50482 46900 50494
rect 46844 50430 46846 50482
rect 46898 50430 46900 50482
rect 46172 49922 46564 49924
rect 46172 49870 46174 49922
rect 46226 49870 46564 49922
rect 46172 49868 46564 49870
rect 46172 49858 46228 49868
rect 46060 49532 46452 49588
rect 46172 49028 46228 49038
rect 46172 48934 46228 48972
rect 45836 48916 45892 48926
rect 45836 48822 45892 48860
rect 46396 48914 46452 49532
rect 46396 48862 46398 48914
rect 46450 48862 46452 48914
rect 46396 48850 46452 48862
rect 46172 48466 46228 48478
rect 46172 48414 46174 48466
rect 46226 48414 46228 48466
rect 46060 48244 46116 48254
rect 46060 48150 46116 48188
rect 46172 47684 46228 48414
rect 46284 48132 46340 48142
rect 46284 47684 46340 48076
rect 46284 47628 46452 47684
rect 46172 47618 46228 47628
rect 45948 47460 46004 47470
rect 45948 47366 46004 47404
rect 46060 47012 46116 47022
rect 45836 46900 45892 46910
rect 45836 46806 45892 46844
rect 46060 46674 46116 46956
rect 46060 46622 46062 46674
rect 46114 46622 46116 46674
rect 46060 45890 46116 46622
rect 46060 45838 46062 45890
rect 46114 45838 46116 45890
rect 46060 45826 46116 45838
rect 45724 45612 45892 45668
rect 45724 45220 45780 45230
rect 45724 45126 45780 45164
rect 45836 44324 45892 45612
rect 45836 44230 45892 44268
rect 46060 44098 46116 44110
rect 46060 44046 46062 44098
rect 46114 44046 46116 44098
rect 46060 43764 46116 44046
rect 46060 43698 46116 43708
rect 46172 43428 46228 43438
rect 46172 43334 46228 43372
rect 45836 42980 45892 42990
rect 45836 42886 45892 42924
rect 45388 42028 45668 42084
rect 44940 39900 45108 39956
rect 45276 41972 45332 41982
rect 45388 41972 45444 42028
rect 45276 41970 45444 41972
rect 45276 41918 45278 41970
rect 45330 41918 45444 41970
rect 45276 41916 45444 41918
rect 45724 41972 45780 41982
rect 45276 40402 45332 41916
rect 45724 41878 45780 41916
rect 45948 41970 46004 41982
rect 45948 41918 45950 41970
rect 46002 41918 46004 41970
rect 45948 41748 46004 41918
rect 46284 41970 46340 41982
rect 46284 41918 46286 41970
rect 46338 41918 46340 41970
rect 46284 41860 46340 41918
rect 46396 41972 46452 47628
rect 46508 42420 46564 49868
rect 46844 49812 46900 50430
rect 46956 50484 47012 50494
rect 47180 50428 47236 51548
rect 47516 51378 47572 51884
rect 47628 51874 47684 51884
rect 47516 51326 47518 51378
rect 47570 51326 47572 51378
rect 47516 51268 47572 51326
rect 47516 50708 47572 51212
rect 47516 50642 47572 50652
rect 47964 51268 48020 51278
rect 48076 51268 48132 53900
rect 49084 53618 49140 53630
rect 49084 53566 49086 53618
rect 49138 53566 49140 53618
rect 48188 52276 48244 52286
rect 48188 52182 48244 52220
rect 49084 52276 49140 53566
rect 49084 52210 49140 52220
rect 48860 52164 48916 52174
rect 47964 51266 48132 51268
rect 47964 51214 47966 51266
rect 48018 51214 48132 51266
rect 47964 51212 48132 51214
rect 48636 51492 48692 51502
rect 48636 51378 48692 51436
rect 48636 51326 48638 51378
rect 48690 51326 48692 51378
rect 47292 50596 47348 50606
rect 47292 50502 47348 50540
rect 47964 50428 48020 51212
rect 48636 50818 48692 51326
rect 48860 51154 48916 52108
rect 49196 51380 49252 51390
rect 48860 51102 48862 51154
rect 48914 51102 48916 51154
rect 48860 51090 48916 51102
rect 49084 51378 49252 51380
rect 49084 51326 49198 51378
rect 49250 51326 49252 51378
rect 49084 51324 49252 51326
rect 48636 50766 48638 50818
rect 48690 50766 48692 50818
rect 48636 50754 48692 50766
rect 46956 50034 47012 50428
rect 46956 49982 46958 50034
rect 47010 49982 47012 50034
rect 46956 49970 47012 49982
rect 47068 50372 47236 50428
rect 47628 50372 48020 50428
rect 48076 50708 48132 50718
rect 48076 50484 48132 50652
rect 48860 50594 48916 50606
rect 48860 50542 48862 50594
rect 48914 50542 48916 50594
rect 48412 50484 48468 50494
rect 48860 50484 48916 50542
rect 49084 50596 49140 51324
rect 49196 51314 49252 51324
rect 49084 50502 49140 50540
rect 48076 50482 48580 50484
rect 48076 50430 48078 50482
rect 48130 50430 48414 50482
rect 48466 50430 48580 50482
rect 48076 50428 48580 50430
rect 48076 50418 48132 50428
rect 48412 50418 48468 50428
rect 46844 49718 46900 49756
rect 46732 48914 46788 48926
rect 46732 48862 46734 48914
rect 46786 48862 46788 48914
rect 46732 48132 46788 48862
rect 47068 48468 47124 50372
rect 47180 49028 47236 49038
rect 47180 48934 47236 48972
rect 47068 48466 47348 48468
rect 47068 48414 47070 48466
rect 47122 48414 47348 48466
rect 47068 48412 47348 48414
rect 47068 48402 47124 48412
rect 46732 48038 46788 48076
rect 46844 48020 46900 48030
rect 46732 47572 46788 47582
rect 46844 47572 46900 47964
rect 46732 47570 46900 47572
rect 46732 47518 46734 47570
rect 46786 47518 46900 47570
rect 46732 47516 46900 47518
rect 46732 47506 46788 47516
rect 46956 47458 47012 47470
rect 46956 47406 46958 47458
rect 47010 47406 47012 47458
rect 46956 47124 47012 47406
rect 47180 47460 47236 47470
rect 47180 47366 47236 47404
rect 46956 47058 47012 47068
rect 47292 45892 47348 48412
rect 47404 48242 47460 48254
rect 47404 48190 47406 48242
rect 47458 48190 47460 48242
rect 47404 48020 47460 48190
rect 47404 47954 47460 47964
rect 47404 47684 47460 47694
rect 47404 47590 47460 47628
rect 47404 45892 47460 45902
rect 47180 45890 47460 45892
rect 47180 45838 47406 45890
rect 47458 45838 47460 45890
rect 47180 45836 47460 45838
rect 46844 45220 46900 45230
rect 46844 45106 46900 45164
rect 46844 45054 46846 45106
rect 46898 45054 46900 45106
rect 46620 44994 46676 45006
rect 46620 44942 46622 44994
rect 46674 44942 46676 44994
rect 46620 44884 46676 44942
rect 46620 44818 46676 44828
rect 46732 44996 46788 45006
rect 46732 44546 46788 44940
rect 46732 44494 46734 44546
rect 46786 44494 46788 44546
rect 46732 44482 46788 44494
rect 46844 44548 46900 45054
rect 47068 45108 47124 45118
rect 47068 45014 47124 45052
rect 47180 44884 47236 45836
rect 47404 45826 47460 45836
rect 47404 45108 47460 45118
rect 46956 44548 47012 44558
rect 46844 44546 47012 44548
rect 46844 44494 46958 44546
rect 47010 44494 47012 44546
rect 46844 44492 47012 44494
rect 46956 44482 47012 44492
rect 47180 44324 47236 44828
rect 47292 44882 47348 44894
rect 47292 44830 47294 44882
rect 47346 44830 47348 44882
rect 47292 44548 47348 44830
rect 47292 44482 47348 44492
rect 47404 44546 47460 45052
rect 47404 44494 47406 44546
rect 47458 44494 47460 44546
rect 47404 44482 47460 44494
rect 47516 44548 47572 44558
rect 47516 44454 47572 44492
rect 47292 44324 47348 44334
rect 47180 44322 47348 44324
rect 47180 44270 47294 44322
rect 47346 44270 47348 44322
rect 47180 44268 47348 44270
rect 47292 44258 47348 44268
rect 46732 43764 46788 43774
rect 46732 43670 46788 43708
rect 46508 42354 46564 42364
rect 46508 42196 46564 42206
rect 46508 42194 46676 42196
rect 46508 42142 46510 42194
rect 46562 42142 46676 42194
rect 46508 42140 46676 42142
rect 46508 42130 46564 42140
rect 46396 41916 46564 41972
rect 46284 41804 46452 41860
rect 45612 41692 46004 41748
rect 46172 41748 46228 41758
rect 45612 41186 45668 41692
rect 46172 41654 46228 41692
rect 46396 41188 46452 41804
rect 45612 41134 45614 41186
rect 45666 41134 45668 41186
rect 45612 40628 45668 41134
rect 45612 40562 45668 40572
rect 45836 41186 46452 41188
rect 45836 41134 46398 41186
rect 46450 41134 46452 41186
rect 45836 41132 46452 41134
rect 45836 40514 45892 41132
rect 46396 41122 46452 41132
rect 45836 40462 45838 40514
rect 45890 40462 45892 40514
rect 45836 40450 45892 40462
rect 46284 40964 46340 40974
rect 45276 40350 45278 40402
rect 45330 40350 45332 40402
rect 44828 39396 44884 39406
rect 44716 39394 44884 39396
rect 44716 39342 44830 39394
rect 44882 39342 44884 39394
rect 44716 39340 44884 39342
rect 44716 38834 44772 39340
rect 44828 39330 44884 39340
rect 44716 38782 44718 38834
rect 44770 38782 44772 38834
rect 44716 38668 44772 38782
rect 43820 38612 44436 38668
rect 44492 38612 44660 38668
rect 44716 38612 44884 38668
rect 43484 38050 43652 38052
rect 43484 37998 43486 38050
rect 43538 37998 43652 38050
rect 43484 37996 43652 37998
rect 43484 37986 43540 37996
rect 43372 35858 43428 35868
rect 43092 35084 43204 35140
rect 43260 35586 43316 35598
rect 43260 35534 43262 35586
rect 43314 35534 43316 35586
rect 41356 35028 41412 35038
rect 41356 34130 41412 34972
rect 41356 34078 41358 34130
rect 41410 34078 41412 34130
rect 41356 34066 41412 34078
rect 42476 33348 42532 33358
rect 42476 33254 42532 33292
rect 43036 33346 43092 35084
rect 43260 34356 43316 35534
rect 43372 34916 43428 34926
rect 43596 34916 43652 37996
rect 44044 37492 44100 37502
rect 43372 34914 43540 34916
rect 43372 34862 43374 34914
rect 43426 34862 43540 34914
rect 43372 34860 43540 34862
rect 43596 34860 43764 34916
rect 43372 34850 43428 34860
rect 43260 34290 43316 34300
rect 43036 33294 43038 33346
rect 43090 33294 43092 33346
rect 43036 33282 43092 33294
rect 43148 33236 43204 33274
rect 43148 33170 43204 33180
rect 43484 33124 43540 34860
rect 43596 34692 43652 34702
rect 43596 34598 43652 34636
rect 43708 34468 43764 34860
rect 43596 34412 43764 34468
rect 43932 34692 43988 34702
rect 43596 33572 43652 34412
rect 43932 34354 43988 34636
rect 43932 34302 43934 34354
rect 43986 34302 43988 34354
rect 43932 33684 43988 34302
rect 43932 33618 43988 33628
rect 43596 33516 43876 33572
rect 43708 33346 43764 33358
rect 43708 33294 43710 33346
rect 43762 33294 43764 33346
rect 43372 33122 43540 33124
rect 43372 33070 43486 33122
rect 43538 33070 43540 33122
rect 43372 33068 43540 33070
rect 43148 33012 43204 33022
rect 43148 32786 43204 32956
rect 43148 32734 43150 32786
rect 43202 32734 43204 32786
rect 43148 32722 43204 32734
rect 42700 32228 42756 32238
rect 41692 31220 41748 31230
rect 41692 31126 41748 31164
rect 41916 31220 41972 31230
rect 41916 31126 41972 31164
rect 41244 31054 41246 31106
rect 41298 31054 41300 31106
rect 41244 31042 41300 31054
rect 39788 30996 39844 31006
rect 39788 30882 39844 30940
rect 41356 30996 41412 31006
rect 41356 30902 41412 30940
rect 42028 30996 42084 31006
rect 42028 30994 42196 30996
rect 42028 30942 42030 30994
rect 42082 30942 42196 30994
rect 42028 30940 42196 30942
rect 42028 30930 42084 30940
rect 40348 30884 40404 30894
rect 39788 30830 39790 30882
rect 39842 30830 39844 30882
rect 39788 30818 39844 30830
rect 40236 30828 40348 30884
rect 39676 30370 39732 30380
rect 38556 30212 38612 30222
rect 37660 29986 38388 29988
rect 37660 29934 37662 29986
rect 37714 29934 38388 29986
rect 37660 29932 38388 29934
rect 37660 29922 37716 29932
rect 37324 29586 37380 29596
rect 38332 29538 38388 29932
rect 38444 30210 38612 30212
rect 38444 30158 38558 30210
rect 38610 30158 38612 30210
rect 38444 30156 38612 30158
rect 38444 29652 38500 30156
rect 38556 30146 38612 30156
rect 40236 30098 40292 30828
rect 40348 30818 40404 30828
rect 41020 30884 41076 30894
rect 41020 30790 41076 30828
rect 42140 30434 42196 30940
rect 42140 30382 42142 30434
rect 42194 30382 42196 30434
rect 42140 30370 42196 30382
rect 42700 30994 42756 32172
rect 42700 30942 42702 30994
rect 42754 30942 42756 30994
rect 40236 30046 40238 30098
rect 40290 30046 40292 30098
rect 40236 30034 40292 30046
rect 38444 29558 38500 29596
rect 38556 29988 38612 29998
rect 38332 29486 38334 29538
rect 38386 29486 38388 29538
rect 33740 29428 33796 29438
rect 33740 29334 33796 29372
rect 37884 29316 37940 29326
rect 37324 29314 37940 29316
rect 37324 29262 37886 29314
rect 37938 29262 37940 29314
rect 37324 29260 37940 29262
rect 36876 29202 36932 29214
rect 36876 29150 36878 29202
rect 36930 29150 36932 29202
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 33964 28756 34020 28766
rect 33964 28662 34020 28700
rect 33516 28590 33518 28642
rect 33570 28590 33572 28642
rect 33516 28578 33572 28590
rect 34972 28644 35028 28654
rect 33180 28478 33182 28530
rect 33234 28478 33236 28530
rect 33180 28466 33236 28478
rect 32956 28420 33012 28430
rect 32956 28326 33012 28364
rect 32620 28030 32622 28082
rect 32674 28030 32676 28082
rect 32620 28018 32676 28030
rect 33964 28084 34020 28094
rect 31276 27022 31278 27074
rect 31330 27022 31332 27074
rect 31276 27010 31332 27022
rect 31724 27188 31780 27198
rect 31724 27074 31780 27132
rect 31724 27022 31726 27074
rect 31778 27022 31780 27074
rect 31724 27010 31780 27022
rect 32284 27188 32340 27198
rect 30716 26962 30772 26974
rect 30716 26910 30718 26962
rect 30770 26910 30772 26962
rect 30716 26908 30772 26910
rect 30604 26852 30772 26908
rect 29148 25620 29204 25630
rect 29148 25508 29204 25564
rect 28588 25414 28644 25452
rect 28812 25506 29204 25508
rect 28812 25454 29150 25506
rect 29202 25454 29204 25506
rect 28812 25452 29204 25454
rect 28252 25106 28308 25116
rect 28364 25396 28420 25406
rect 28364 24834 28420 25340
rect 28364 24782 28366 24834
rect 28418 24782 28420 24834
rect 28140 24050 28196 24062
rect 28140 23998 28142 24050
rect 28194 23998 28196 24050
rect 28140 23156 28196 23998
rect 28364 23268 28420 24782
rect 28476 25172 28532 25182
rect 28476 23938 28532 25116
rect 28700 24836 28756 24846
rect 28700 24742 28756 24780
rect 28476 23886 28478 23938
rect 28530 23886 28532 23938
rect 28476 23874 28532 23886
rect 28420 23212 28532 23268
rect 28364 23202 28420 23212
rect 28252 23156 28308 23166
rect 28196 23154 28308 23156
rect 28196 23102 28254 23154
rect 28306 23102 28308 23154
rect 28196 23100 28308 23102
rect 28140 23062 28196 23100
rect 28252 23090 28308 23100
rect 28028 22876 28420 22932
rect 28028 22260 28084 22270
rect 28028 22258 28308 22260
rect 28028 22206 28030 22258
rect 28082 22206 28308 22258
rect 28028 22204 28308 22206
rect 28028 22194 28084 22204
rect 27916 21980 28196 22036
rect 27804 21758 27806 21810
rect 27858 21758 27860 21810
rect 27804 21746 27860 21758
rect 28028 20804 28084 20814
rect 27692 20626 27748 20636
rect 27804 20802 28084 20804
rect 27804 20750 28030 20802
rect 28082 20750 28084 20802
rect 27804 20748 28084 20750
rect 27580 20356 27636 20366
rect 27580 20188 27636 20300
rect 27580 20132 27748 20188
rect 27468 20038 27524 20076
rect 27580 20018 27636 20030
rect 27580 19966 27582 20018
rect 27634 19966 27636 20018
rect 27580 19908 27636 19966
rect 27580 19572 27636 19852
rect 27468 19516 27636 19572
rect 27692 20018 27748 20132
rect 27692 19966 27694 20018
rect 27746 19966 27748 20018
rect 27468 18900 27524 19516
rect 27580 19348 27636 19358
rect 27692 19348 27748 19966
rect 27580 19346 27748 19348
rect 27580 19294 27582 19346
rect 27634 19294 27748 19346
rect 27580 19292 27748 19294
rect 27580 19282 27636 19292
rect 27468 18834 27524 18844
rect 27692 18564 27748 18574
rect 27692 18340 27748 18508
rect 27692 18246 27748 18284
rect 27692 17332 27748 17342
rect 27580 16994 27636 17006
rect 27580 16942 27582 16994
rect 27634 16942 27636 16994
rect 27244 12684 27412 12740
rect 27468 16772 27524 16782
rect 27244 11732 27300 12684
rect 27356 12516 27412 12526
rect 27356 12402 27412 12460
rect 27356 12350 27358 12402
rect 27410 12350 27412 12402
rect 27356 12068 27412 12350
rect 27356 12002 27412 12012
rect 27468 11844 27524 16716
rect 27580 16212 27636 16942
rect 27580 16146 27636 16156
rect 27692 16884 27748 17276
rect 27804 17220 27860 20748
rect 28028 20738 28084 20748
rect 28140 20580 28196 21980
rect 28028 20524 28196 20580
rect 28028 20188 28084 20524
rect 27804 17154 27860 17164
rect 27916 20132 28084 20188
rect 28140 20132 28196 20142
rect 27804 16884 27860 16894
rect 27692 16882 27860 16884
rect 27692 16830 27806 16882
rect 27858 16830 27860 16882
rect 27692 16828 27860 16830
rect 27580 15986 27636 15998
rect 27580 15934 27582 15986
rect 27634 15934 27636 15986
rect 27580 15428 27636 15934
rect 27692 15876 27748 16828
rect 27804 16818 27860 16828
rect 27916 16772 27972 20132
rect 28140 20038 28196 20076
rect 28140 19572 28196 19582
rect 28252 19572 28308 22204
rect 28364 21812 28420 22876
rect 28476 22370 28532 23212
rect 28476 22318 28478 22370
rect 28530 22318 28532 22370
rect 28476 22306 28532 22318
rect 28364 21810 28644 21812
rect 28364 21758 28366 21810
rect 28418 21758 28644 21810
rect 28364 21756 28644 21758
rect 28364 20356 28420 21756
rect 28588 21586 28644 21756
rect 28588 21534 28590 21586
rect 28642 21534 28644 21586
rect 28588 21522 28644 21534
rect 28476 20804 28532 20814
rect 28476 20710 28532 20748
rect 28364 20290 28420 20300
rect 28812 20188 28868 25452
rect 29148 25442 29204 25452
rect 29260 25396 29316 25406
rect 29260 25302 29316 25340
rect 29260 24948 29316 24958
rect 29372 24948 29428 26236
rect 30380 26292 30436 26302
rect 30380 26198 30436 26236
rect 30268 25956 30324 25966
rect 29708 25844 29764 25854
rect 29260 24946 29428 24948
rect 29260 24894 29262 24946
rect 29314 24894 29428 24946
rect 29260 24892 29428 24894
rect 29596 25172 29652 25182
rect 29260 24882 29316 24892
rect 29148 23938 29204 23950
rect 29148 23886 29150 23938
rect 29202 23886 29204 23938
rect 29036 23042 29092 23054
rect 29036 22990 29038 23042
rect 29090 22990 29092 23042
rect 28588 20132 28644 20142
rect 28588 20038 28644 20076
rect 28700 20132 28868 20188
rect 28924 21698 28980 21710
rect 28924 21646 28926 21698
rect 28978 21646 28980 21698
rect 28196 19516 28308 19572
rect 28140 19346 28196 19516
rect 28140 19294 28142 19346
rect 28194 19294 28196 19346
rect 28140 19282 28196 19294
rect 28476 19236 28532 19246
rect 28476 18674 28532 19180
rect 28588 19010 28644 19022
rect 28588 18958 28590 19010
rect 28642 18958 28644 19010
rect 28588 18788 28644 18958
rect 28588 18722 28644 18732
rect 28476 18622 28478 18674
rect 28530 18622 28532 18674
rect 28476 18610 28532 18622
rect 28028 18338 28084 18350
rect 28028 18286 28030 18338
rect 28082 18286 28084 18338
rect 28028 16996 28084 18286
rect 28252 17892 28308 17902
rect 28252 17798 28308 17836
rect 28028 16930 28084 16940
rect 28364 17220 28420 17230
rect 27916 16716 28084 16772
rect 27916 16212 27972 16222
rect 27804 16100 27860 16110
rect 27804 16006 27860 16044
rect 27692 15820 27860 15876
rect 27580 15362 27636 15372
rect 27692 15652 27748 15662
rect 27692 15426 27748 15596
rect 27692 15374 27694 15426
rect 27746 15374 27748 15426
rect 27692 15362 27748 15374
rect 27804 14644 27860 15820
rect 27692 14588 27860 14644
rect 27916 15316 27972 16156
rect 27692 13412 27748 14588
rect 27804 14420 27860 14430
rect 27804 14326 27860 14364
rect 27244 11666 27300 11676
rect 27356 11788 27524 11844
rect 27580 12962 27636 12974
rect 27580 12910 27582 12962
rect 27634 12910 27636 12962
rect 27580 12292 27636 12910
rect 27692 12964 27748 13356
rect 27692 12898 27748 12908
rect 27804 13748 27860 13758
rect 27916 13748 27972 15260
rect 27860 13692 27972 13748
rect 28028 14642 28084 16716
rect 28140 15540 28196 15578
rect 28140 15474 28196 15484
rect 28364 15428 28420 17164
rect 28700 17108 28756 20132
rect 28812 20018 28868 20030
rect 28812 19966 28814 20018
rect 28866 19966 28868 20018
rect 28812 18452 28868 19966
rect 28924 19908 28980 21646
rect 28924 19842 28980 19852
rect 28812 18386 28868 18396
rect 28252 15372 28420 15428
rect 28588 17052 28756 17108
rect 28588 15652 28644 17052
rect 28700 16882 28756 16894
rect 28700 16830 28702 16882
rect 28754 16830 28756 16882
rect 28700 16548 28756 16830
rect 28700 16482 28756 16492
rect 29036 16212 29092 22990
rect 29148 22594 29204 23886
rect 29596 23938 29652 25116
rect 29596 23886 29598 23938
rect 29650 23886 29652 23938
rect 29596 23874 29652 23886
rect 29708 24946 29764 25788
rect 29708 24894 29710 24946
rect 29762 24894 29764 24946
rect 29484 23268 29540 23278
rect 29484 23174 29540 23212
rect 29148 22542 29150 22594
rect 29202 22542 29204 22594
rect 29148 22530 29204 22542
rect 29260 22260 29316 22270
rect 29260 22166 29316 22204
rect 29596 21810 29652 21822
rect 29596 21758 29598 21810
rect 29650 21758 29652 21810
rect 29148 21698 29204 21710
rect 29148 21646 29150 21698
rect 29202 21646 29204 21698
rect 29148 21476 29204 21646
rect 29148 20916 29204 21420
rect 29148 20850 29204 20860
rect 29596 20802 29652 21758
rect 29596 20750 29598 20802
rect 29650 20750 29652 20802
rect 29596 20738 29652 20750
rect 29708 20188 29764 24894
rect 29932 25620 29988 25630
rect 29932 24612 29988 25564
rect 30044 25508 30100 25518
rect 30044 25414 30100 25452
rect 30156 25282 30212 25294
rect 30156 25230 30158 25282
rect 30210 25230 30212 25282
rect 30156 24836 30212 25230
rect 30156 24770 30212 24780
rect 30156 24612 30212 24622
rect 29932 24610 30212 24612
rect 29932 24558 30158 24610
rect 30210 24558 30212 24610
rect 29932 24556 30212 24558
rect 30156 24546 30212 24556
rect 29932 23154 29988 23166
rect 29932 23102 29934 23154
rect 29986 23102 29988 23154
rect 29932 22596 29988 23102
rect 29932 22530 29988 22540
rect 29820 22482 29876 22494
rect 29820 22430 29822 22482
rect 29874 22430 29876 22482
rect 29820 22370 29876 22430
rect 29820 22318 29822 22370
rect 29874 22318 29876 22370
rect 29820 21700 29876 22318
rect 29820 20804 29876 21644
rect 29820 20738 29876 20748
rect 30044 21586 30100 21598
rect 30044 21534 30046 21586
rect 30098 21534 30100 21586
rect 29708 20132 29876 20188
rect 29148 19572 29204 19582
rect 29148 18450 29204 19516
rect 29148 18398 29150 18450
rect 29202 18398 29204 18450
rect 29148 18386 29204 18398
rect 29260 19234 29316 19246
rect 29596 19236 29652 19246
rect 29260 19182 29262 19234
rect 29314 19182 29316 19234
rect 29260 18788 29316 19182
rect 29484 19234 29652 19236
rect 29484 19182 29598 19234
rect 29650 19182 29652 19234
rect 29484 19180 29652 19182
rect 29484 18900 29540 19180
rect 29596 19170 29652 19180
rect 29260 17220 29316 18732
rect 29372 18844 29540 18900
rect 29596 19010 29652 19022
rect 29596 18958 29598 19010
rect 29650 18958 29652 19010
rect 29372 18450 29428 18844
rect 29484 18676 29540 18686
rect 29484 18562 29540 18620
rect 29484 18510 29486 18562
rect 29538 18510 29540 18562
rect 29484 18498 29540 18510
rect 29372 18398 29374 18450
rect 29426 18398 29428 18450
rect 29372 17444 29428 18398
rect 29484 17668 29540 17678
rect 29596 17668 29652 18958
rect 29820 18452 29876 20132
rect 30044 20020 30100 21534
rect 30044 19954 30100 19964
rect 29932 19572 29988 19582
rect 29932 19234 29988 19516
rect 29932 19182 29934 19234
rect 29986 19182 29988 19234
rect 29932 19170 29988 19182
rect 29820 18396 30100 18452
rect 29932 18226 29988 18238
rect 29932 18174 29934 18226
rect 29986 18174 29988 18226
rect 29484 17666 29652 17668
rect 29484 17614 29486 17666
rect 29538 17614 29652 17666
rect 29484 17612 29652 17614
rect 29708 17780 29764 17790
rect 29484 17602 29540 17612
rect 29372 17388 29540 17444
rect 28140 15314 28196 15326
rect 28140 15262 28142 15314
rect 28194 15262 28196 15314
rect 28140 14980 28196 15262
rect 28140 14914 28196 14924
rect 28028 14590 28030 14642
rect 28082 14590 28084 14642
rect 27132 10670 27134 10722
rect 27186 10670 27188 10722
rect 27132 10658 27188 10670
rect 27244 11508 27300 11518
rect 27020 10558 27022 10610
rect 27074 10558 27076 10610
rect 27020 10546 27076 10558
rect 26908 10500 26964 10510
rect 26908 9828 26964 10444
rect 27244 10164 27300 11452
rect 27356 11394 27412 11788
rect 27580 11620 27636 12236
rect 27692 12740 27748 12750
rect 27692 12290 27748 12684
rect 27804 12402 27860 13692
rect 27804 12350 27806 12402
rect 27858 12350 27860 12402
rect 27804 12338 27860 12350
rect 27916 13076 27972 13086
rect 27692 12238 27694 12290
rect 27746 12238 27748 12290
rect 27692 12226 27748 12238
rect 27804 12180 27860 12190
rect 27804 11954 27860 12124
rect 27804 11902 27806 11954
rect 27858 11902 27860 11954
rect 27804 11890 27860 11902
rect 27356 11342 27358 11394
rect 27410 11342 27412 11394
rect 27356 11330 27412 11342
rect 27468 11564 27636 11620
rect 27468 11172 27524 11564
rect 27916 11282 27972 13020
rect 27916 11230 27918 11282
rect 27970 11230 27972 11282
rect 27916 11218 27972 11230
rect 27132 10108 27300 10164
rect 27356 11116 27524 11172
rect 27580 11172 27636 11182
rect 27020 9828 27076 9838
rect 26908 9826 27076 9828
rect 26908 9774 27022 9826
rect 27074 9774 27076 9826
rect 26908 9772 27076 9774
rect 27020 9762 27076 9772
rect 26796 9660 26964 9716
rect 26796 9268 26852 9278
rect 26796 9174 26852 9212
rect 26684 8754 26740 8764
rect 26796 8708 26852 8718
rect 26796 6916 26852 8652
rect 26572 6850 26628 6860
rect 26684 6860 26852 6916
rect 26908 8260 26964 9660
rect 27132 9266 27188 10108
rect 27356 10052 27412 11116
rect 27580 11078 27636 11116
rect 27244 9996 27412 10052
rect 27580 10052 27636 10062
rect 27244 9826 27300 9996
rect 27244 9774 27246 9826
rect 27298 9774 27300 9826
rect 27244 9762 27300 9774
rect 27468 9940 27524 9950
rect 27468 9826 27524 9884
rect 27468 9774 27470 9826
rect 27522 9774 27524 9826
rect 27468 9762 27524 9774
rect 27356 9602 27412 9614
rect 27356 9550 27358 9602
rect 27410 9550 27412 9602
rect 27356 9380 27412 9550
rect 27356 9314 27412 9324
rect 27132 9214 27134 9266
rect 27186 9214 27188 9266
rect 27132 9202 27188 9214
rect 27580 9266 27636 9996
rect 28028 9940 28084 14590
rect 28140 14308 28196 14318
rect 28140 13858 28196 14252
rect 28140 13806 28142 13858
rect 28194 13806 28196 13858
rect 28140 13794 28196 13806
rect 28140 12964 28196 12974
rect 28140 12628 28196 12908
rect 28140 12562 28196 12572
rect 28252 12404 28308 15372
rect 28364 15204 28420 15214
rect 28364 15092 28532 15148
rect 28476 14530 28532 15092
rect 28476 14478 28478 14530
rect 28530 14478 28532 14530
rect 28476 14466 28532 14478
rect 28588 13972 28644 15596
rect 28700 16156 29092 16212
rect 29148 17164 29316 17220
rect 28700 15314 28756 16156
rect 28700 15262 28702 15314
rect 28754 15262 28756 15314
rect 28700 15148 28756 15262
rect 28924 15988 28980 15998
rect 28924 15314 28980 15932
rect 28924 15262 28926 15314
rect 28978 15262 28980 15314
rect 28924 15250 28980 15262
rect 29036 15876 29092 15886
rect 28700 15092 28868 15148
rect 28588 13916 28756 13972
rect 28476 13746 28532 13758
rect 28476 13694 28478 13746
rect 28530 13694 28532 13746
rect 28476 13188 28532 13694
rect 28588 13636 28644 13646
rect 28588 13542 28644 13580
rect 28476 13122 28532 13132
rect 28700 13074 28756 13916
rect 28812 13412 28868 15092
rect 28924 13412 28980 13422
rect 28812 13356 28924 13412
rect 28700 13022 28702 13074
rect 28754 13022 28756 13074
rect 28700 13010 28756 13022
rect 28140 12402 28308 12404
rect 28140 12350 28254 12402
rect 28306 12350 28308 12402
rect 28140 12348 28308 12350
rect 28140 10610 28196 12348
rect 28252 12338 28308 12348
rect 28700 12066 28756 12078
rect 28700 12014 28702 12066
rect 28754 12014 28756 12066
rect 28700 11956 28756 12014
rect 28700 11890 28756 11900
rect 28812 11844 28868 11854
rect 28924 11844 28980 13356
rect 28868 11788 28980 11844
rect 28140 10558 28142 10610
rect 28194 10558 28196 10610
rect 28140 10546 28196 10558
rect 28476 11732 28532 11742
rect 27804 9884 28084 9940
rect 28476 9938 28532 11676
rect 28700 11508 28756 11518
rect 28588 11452 28700 11508
rect 28588 11394 28644 11452
rect 28588 11342 28590 11394
rect 28642 11342 28644 11394
rect 28588 11330 28644 11342
rect 28476 9886 28478 9938
rect 28530 9886 28532 9938
rect 27692 9828 27748 9838
rect 27692 9734 27748 9772
rect 27580 9214 27582 9266
rect 27634 9214 27636 9266
rect 27580 9202 27636 9214
rect 27804 8932 27860 9884
rect 28476 9874 28532 9886
rect 28364 9828 28420 9838
rect 28252 9772 28364 9828
rect 27916 9268 27972 9278
rect 27916 9174 27972 9212
rect 28252 9268 28308 9772
rect 28364 9762 28420 9772
rect 28700 9268 28756 11452
rect 28812 11396 28868 11788
rect 28812 10834 28868 11340
rect 28812 10782 28814 10834
rect 28866 10782 28868 10834
rect 28812 10770 28868 10782
rect 29036 10388 29092 15820
rect 29148 13860 29204 17164
rect 29260 16996 29316 17006
rect 29260 16994 29428 16996
rect 29260 16942 29262 16994
rect 29314 16942 29428 16994
rect 29260 16940 29428 16942
rect 29260 16930 29316 16940
rect 29260 16548 29316 16558
rect 29260 16098 29316 16492
rect 29260 16046 29262 16098
rect 29314 16046 29316 16098
rect 29260 15538 29316 16046
rect 29260 15486 29262 15538
rect 29314 15486 29316 15538
rect 29260 15474 29316 15486
rect 29372 15874 29428 16940
rect 29484 15988 29540 17388
rect 29708 17442 29764 17724
rect 29932 17666 29988 18174
rect 29932 17614 29934 17666
rect 29986 17614 29988 17666
rect 29932 17602 29988 17614
rect 29708 17390 29710 17442
rect 29762 17390 29764 17442
rect 29708 17378 29764 17390
rect 29820 17554 29876 17566
rect 29820 17502 29822 17554
rect 29874 17502 29876 17554
rect 29708 16772 29764 16782
rect 29820 16772 29876 17502
rect 29764 16716 29876 16772
rect 29708 16706 29764 16716
rect 29708 16212 29764 16222
rect 29708 16118 29764 16156
rect 29484 15922 29540 15932
rect 29820 16098 29876 16110
rect 29820 16046 29822 16098
rect 29874 16046 29876 16098
rect 29372 15822 29374 15874
rect 29426 15822 29428 15874
rect 29372 15540 29428 15822
rect 29372 15474 29428 15484
rect 29596 15874 29652 15886
rect 29596 15822 29598 15874
rect 29650 15822 29652 15874
rect 29596 15316 29652 15822
rect 29596 15222 29652 15260
rect 29820 15876 29876 16046
rect 29820 15204 29876 15820
rect 29820 15202 29988 15204
rect 29820 15150 29822 15202
rect 29874 15150 29988 15202
rect 29820 15148 29988 15150
rect 29820 15138 29876 15148
rect 29372 14420 29428 14430
rect 29148 13804 29316 13860
rect 29148 13636 29204 13646
rect 29148 10500 29204 13580
rect 29260 12292 29316 13804
rect 29372 13748 29428 14364
rect 29484 14308 29540 14318
rect 29484 14306 29652 14308
rect 29484 14254 29486 14306
rect 29538 14254 29652 14306
rect 29484 14252 29652 14254
rect 29484 14242 29540 14252
rect 29372 12962 29428 13692
rect 29372 12910 29374 12962
rect 29426 12910 29428 12962
rect 29372 12898 29428 12910
rect 29484 13860 29540 13870
rect 29484 12850 29540 13804
rect 29596 13524 29652 14252
rect 29932 13636 29988 15148
rect 29932 13570 29988 13580
rect 29596 13458 29652 13468
rect 30044 13412 30100 18396
rect 30268 17892 30324 25900
rect 30492 25730 30548 25742
rect 30492 25678 30494 25730
rect 30546 25678 30548 25730
rect 30380 19572 30436 19582
rect 30380 19010 30436 19516
rect 30380 18958 30382 19010
rect 30434 18958 30436 19010
rect 30380 18450 30436 18958
rect 30492 18564 30548 25678
rect 30604 25172 30660 26852
rect 31052 26290 31108 26302
rect 31052 26238 31054 26290
rect 31106 26238 31108 26290
rect 30716 26068 30772 26078
rect 30716 25618 30772 26012
rect 31052 26068 31108 26238
rect 31052 26002 31108 26012
rect 31276 26290 31332 26302
rect 31276 26238 31278 26290
rect 31330 26238 31332 26290
rect 31276 25956 31332 26238
rect 31612 26068 31668 26078
rect 31612 26066 31780 26068
rect 31612 26014 31614 26066
rect 31666 26014 31780 26066
rect 31612 26012 31780 26014
rect 31612 26002 31668 26012
rect 31276 25890 31332 25900
rect 30716 25566 30718 25618
rect 30770 25566 30772 25618
rect 30716 25554 30772 25566
rect 31276 25730 31332 25742
rect 31276 25678 31278 25730
rect 31330 25678 31332 25730
rect 31276 25620 31332 25678
rect 31612 25620 31668 25630
rect 31276 25618 31668 25620
rect 31276 25566 31278 25618
rect 31330 25566 31614 25618
rect 31666 25566 31668 25618
rect 31276 25564 31668 25566
rect 31276 25554 31332 25564
rect 31612 25554 31668 25564
rect 31724 25508 31780 26012
rect 32060 25732 32116 25742
rect 31836 25508 31892 25518
rect 31724 25506 31892 25508
rect 31724 25454 31838 25506
rect 31890 25454 31892 25506
rect 31724 25452 31892 25454
rect 31836 25284 31892 25452
rect 31836 25218 31892 25228
rect 30604 25106 30660 25116
rect 30604 24948 30660 24958
rect 30660 24892 30996 24948
rect 30604 24854 30660 24892
rect 30940 24724 30996 24892
rect 31164 24836 31220 24846
rect 31164 24724 31220 24780
rect 31836 24724 31892 24734
rect 30940 24722 31108 24724
rect 30940 24670 30942 24722
rect 30994 24670 31108 24722
rect 30940 24668 31108 24670
rect 30940 24658 30996 24668
rect 31052 24052 31108 24668
rect 31164 24722 31332 24724
rect 31164 24670 31166 24722
rect 31218 24670 31332 24722
rect 31164 24668 31332 24670
rect 31164 24658 31220 24668
rect 31164 24052 31220 24062
rect 31052 23996 31164 24052
rect 31164 23958 31220 23996
rect 31276 23940 31332 24668
rect 31836 24630 31892 24668
rect 31388 24500 31444 24510
rect 31388 24498 31556 24500
rect 31388 24446 31390 24498
rect 31442 24446 31556 24498
rect 31388 24444 31556 24446
rect 31388 24434 31444 24444
rect 31388 23940 31444 23950
rect 31276 23938 31444 23940
rect 31276 23886 31390 23938
rect 31442 23886 31444 23938
rect 31276 23884 31444 23886
rect 31388 23874 31444 23884
rect 31500 23826 31556 24444
rect 31500 23774 31502 23826
rect 31554 23774 31556 23826
rect 31388 23604 31444 23614
rect 31500 23604 31556 23774
rect 31444 23548 31556 23604
rect 31948 23716 32004 23726
rect 31388 23538 31444 23548
rect 31388 23266 31444 23278
rect 31388 23214 31390 23266
rect 31442 23214 31444 23266
rect 30940 23154 30996 23166
rect 30940 23102 30942 23154
rect 30994 23102 30996 23154
rect 30940 22258 30996 23102
rect 31276 23156 31332 23166
rect 31276 23062 31332 23100
rect 30940 22206 30942 22258
rect 30994 22206 30996 22258
rect 30828 21586 30884 21598
rect 30828 21534 30830 21586
rect 30882 21534 30884 21586
rect 30604 21476 30660 21486
rect 30604 21382 30660 21420
rect 30716 20804 30772 20814
rect 30492 18470 30548 18508
rect 30604 20802 30772 20804
rect 30604 20750 30718 20802
rect 30770 20750 30772 20802
rect 30604 20748 30772 20750
rect 30380 18398 30382 18450
rect 30434 18398 30436 18450
rect 30380 18386 30436 18398
rect 30604 18228 30660 20748
rect 30716 20738 30772 20748
rect 30716 20244 30772 20282
rect 30716 20178 30772 20188
rect 30828 20018 30884 21534
rect 30940 20804 30996 22206
rect 31164 21812 31220 21822
rect 31052 21700 31108 21710
rect 31052 21606 31108 21644
rect 31164 21698 31220 21756
rect 31388 21812 31444 23214
rect 31948 23154 32004 23660
rect 31948 23102 31950 23154
rect 32002 23102 32004 23154
rect 31500 22484 31556 22494
rect 31500 22390 31556 22428
rect 31948 22370 32004 23102
rect 32060 23156 32116 25676
rect 32172 25620 32228 25630
rect 32172 25526 32228 25564
rect 32060 23090 32116 23100
rect 31948 22318 31950 22370
rect 32002 22318 32004 22370
rect 31948 22306 32004 22318
rect 32284 22036 32340 27132
rect 33964 26962 34020 28028
rect 33964 26910 33966 26962
rect 34018 26910 34020 26962
rect 33964 26898 34020 26910
rect 34972 27076 35028 28588
rect 35644 28644 35700 28654
rect 35532 28532 35588 28542
rect 35532 28082 35588 28476
rect 35532 28030 35534 28082
rect 35586 28030 35588 28082
rect 35532 28018 35588 28030
rect 35644 27970 35700 28588
rect 35644 27918 35646 27970
rect 35698 27918 35700 27970
rect 35644 27906 35700 27918
rect 36428 27970 36484 27982
rect 36428 27918 36430 27970
rect 36482 27918 36484 27970
rect 35532 27636 35588 27646
rect 35532 27542 35588 27580
rect 35756 27524 35812 27534
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35756 27188 35812 27468
rect 35756 27094 35812 27132
rect 36428 27188 36484 27918
rect 36876 27972 36932 29150
rect 37324 28756 37380 29260
rect 37884 29250 37940 29260
rect 37212 28644 37268 28654
rect 37212 28550 37268 28588
rect 37324 28642 37380 28700
rect 37324 28590 37326 28642
rect 37378 28590 37380 28642
rect 37100 28532 37156 28542
rect 37100 28438 37156 28476
rect 36876 27906 36932 27916
rect 36428 27122 36484 27132
rect 37100 27188 37156 27198
rect 37100 27094 37156 27132
rect 34972 26962 35028 27020
rect 34972 26910 34974 26962
rect 35026 26910 35028 26962
rect 34972 26898 35028 26910
rect 35196 27074 35252 27086
rect 35196 27022 35198 27074
rect 35250 27022 35252 27074
rect 35196 26908 35252 27022
rect 36988 27076 37044 27086
rect 36988 26982 37044 27020
rect 34748 26852 34804 26862
rect 34412 26850 34804 26852
rect 34412 26798 34750 26850
rect 34802 26798 34804 26850
rect 34412 26796 34804 26798
rect 34412 25506 34468 26796
rect 34748 26786 34804 26796
rect 35084 26852 35252 26908
rect 37212 26852 37268 26862
rect 35084 25732 35140 26852
rect 37100 26850 37268 26852
rect 37100 26798 37214 26850
rect 37266 26798 37268 26850
rect 37100 26796 37268 26798
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35084 25676 35252 25732
rect 35196 25620 35252 25676
rect 35196 25554 35252 25564
rect 36092 25620 36148 25630
rect 36092 25526 36148 25564
rect 34412 25454 34414 25506
rect 34466 25454 34468 25506
rect 34076 25284 34132 25294
rect 33964 25282 34132 25284
rect 33964 25230 34078 25282
rect 34130 25230 34132 25282
rect 33964 25228 34132 25230
rect 33404 24836 33460 24846
rect 33404 24834 33572 24836
rect 33404 24782 33406 24834
rect 33458 24782 33572 24834
rect 33404 24780 33572 24782
rect 33404 24770 33460 24780
rect 33180 24724 33236 24734
rect 33180 24630 33236 24668
rect 33404 23940 33460 23950
rect 33516 23940 33572 24780
rect 33852 24724 33908 24734
rect 33740 23940 33796 23950
rect 33516 23884 33740 23940
rect 33404 23846 33460 23884
rect 33740 23266 33796 23884
rect 33740 23214 33742 23266
rect 33794 23214 33796 23266
rect 33740 23202 33796 23214
rect 32508 23156 32564 23166
rect 32508 23062 32564 23100
rect 33516 23154 33572 23166
rect 33516 23102 33518 23154
rect 33570 23102 33572 23154
rect 33516 23044 33572 23102
rect 33628 23156 33684 23166
rect 33628 23062 33684 23100
rect 33068 22932 33124 22942
rect 32956 22930 33124 22932
rect 32956 22878 33070 22930
rect 33122 22878 33124 22930
rect 32956 22876 33124 22878
rect 32396 22484 32452 22494
rect 32396 22258 32452 22428
rect 32396 22206 32398 22258
rect 32450 22206 32452 22258
rect 32396 22194 32452 22206
rect 31388 21746 31444 21756
rect 32060 21980 32340 22036
rect 32060 21810 32116 21980
rect 32060 21758 32062 21810
rect 32114 21758 32116 21810
rect 32060 21746 32116 21758
rect 32172 21812 32228 21822
rect 31164 21646 31166 21698
rect 31218 21646 31220 21698
rect 31164 21252 31220 21646
rect 31724 21476 31780 21486
rect 31164 21186 31220 21196
rect 31500 21474 31780 21476
rect 31500 21422 31726 21474
rect 31778 21422 31780 21474
rect 31500 21420 31780 21422
rect 30940 20738 30996 20748
rect 31052 20692 31108 20702
rect 31052 20188 31108 20636
rect 30828 19966 30830 20018
rect 30882 19966 30884 20018
rect 30828 19954 30884 19966
rect 30940 20132 31108 20188
rect 31500 20188 31556 21420
rect 31724 21410 31780 21420
rect 31612 21252 31668 21262
rect 31612 20802 31668 21196
rect 31836 21028 31892 21038
rect 31612 20750 31614 20802
rect 31666 20750 31668 20802
rect 31612 20738 31668 20750
rect 31724 21026 31892 21028
rect 31724 20974 31838 21026
rect 31890 20974 31892 21026
rect 31724 20972 31892 20974
rect 31724 20244 31780 20972
rect 31836 20962 31892 20972
rect 32172 20916 32228 21756
rect 32284 21700 32340 21980
rect 32396 21700 32452 21710
rect 32284 21698 32452 21700
rect 32284 21646 32398 21698
rect 32450 21646 32452 21698
rect 32284 21644 32452 21646
rect 32396 21028 32452 21644
rect 32508 21364 32564 21374
rect 32508 21270 32564 21308
rect 32396 20962 32452 20972
rect 32060 20860 32228 20916
rect 31948 20804 32004 20814
rect 31948 20690 32004 20748
rect 31948 20638 31950 20690
rect 32002 20638 32004 20690
rect 31948 20626 32004 20638
rect 31500 20132 31668 20188
rect 31724 20178 31780 20188
rect 31836 20244 31892 20254
rect 32060 20244 32116 20860
rect 32284 20804 32340 20814
rect 31836 20242 32116 20244
rect 31836 20190 31838 20242
rect 31890 20190 32116 20242
rect 31836 20188 32116 20190
rect 32172 20468 32228 20478
rect 31836 20178 31892 20188
rect 30940 19460 30996 20132
rect 30604 18162 30660 18172
rect 30828 19404 30996 19460
rect 31612 20018 31668 20132
rect 31612 19966 31614 20018
rect 31666 19966 31668 20018
rect 30268 17836 30660 17892
rect 30380 17666 30436 17678
rect 30380 17614 30382 17666
rect 30434 17614 30436 17666
rect 30268 16882 30324 16894
rect 30268 16830 30270 16882
rect 30322 16830 30324 16882
rect 30268 16100 30324 16830
rect 30380 16212 30436 17614
rect 30380 16146 30436 16156
rect 30492 16996 30548 17006
rect 30156 16044 30324 16100
rect 30156 15538 30212 16044
rect 30268 15876 30324 15886
rect 30492 15876 30548 16940
rect 30268 15874 30548 15876
rect 30268 15822 30270 15874
rect 30322 15822 30548 15874
rect 30268 15820 30548 15822
rect 30268 15810 30324 15820
rect 30156 15486 30158 15538
rect 30210 15486 30212 15538
rect 30156 15474 30212 15486
rect 30492 15092 30548 15102
rect 30492 14418 30548 15036
rect 30492 14366 30494 14418
rect 30546 14366 30548 14418
rect 30492 14308 30548 14366
rect 30492 14242 30548 14252
rect 30492 14084 30548 14094
rect 30380 14028 30492 14084
rect 30604 14084 30660 17836
rect 30828 16100 30884 19404
rect 31276 19348 31332 19358
rect 30940 19236 30996 19246
rect 30940 17106 30996 19180
rect 31164 19012 31220 19022
rect 31276 19012 31332 19292
rect 31612 19348 31668 19966
rect 31948 20018 32004 20030
rect 31948 19966 31950 20018
rect 32002 19966 32004 20018
rect 31948 19684 32004 19966
rect 32172 20018 32228 20412
rect 32284 20188 32340 20748
rect 32284 20132 32676 20188
rect 32172 19966 32174 20018
rect 32226 19966 32228 20018
rect 32172 19954 32228 19966
rect 31948 19618 32004 19628
rect 31612 19282 31668 19292
rect 31164 19010 31332 19012
rect 31164 18958 31166 19010
rect 31218 18958 31332 19010
rect 31164 18956 31332 18958
rect 31164 18946 31220 18956
rect 31164 18226 31220 18238
rect 31164 18174 31166 18226
rect 31218 18174 31220 18226
rect 30940 17054 30942 17106
rect 30994 17054 30996 17106
rect 30940 17042 30996 17054
rect 31052 17666 31108 17678
rect 31052 17614 31054 17666
rect 31106 17614 31108 17666
rect 31052 16996 31108 17614
rect 31052 16930 31108 16940
rect 31164 16884 31220 18174
rect 31276 17556 31332 18956
rect 31612 19012 31668 19022
rect 31612 18918 31668 18956
rect 31500 18226 31556 18238
rect 31500 18174 31502 18226
rect 31554 18174 31556 18226
rect 31500 17778 31556 18174
rect 32620 18228 32676 20132
rect 32732 19348 32788 19358
rect 32732 19254 32788 19292
rect 32620 18172 32788 18228
rect 31500 17726 31502 17778
rect 31554 17726 31556 17778
rect 31500 17714 31556 17726
rect 32620 17780 32676 17790
rect 32620 17686 32676 17724
rect 32172 17666 32228 17678
rect 32172 17614 32174 17666
rect 32226 17614 32228 17666
rect 31724 17556 31780 17566
rect 31276 17500 31556 17556
rect 31164 16818 31220 16828
rect 30828 16044 31444 16100
rect 30828 15876 30884 15886
rect 31164 15876 31220 15886
rect 30884 15874 31220 15876
rect 30884 15822 31166 15874
rect 31218 15822 31220 15874
rect 30884 15820 31220 15822
rect 30828 15782 30884 15820
rect 31164 15810 31220 15820
rect 31164 15314 31220 15326
rect 31164 15262 31166 15314
rect 31218 15262 31220 15314
rect 30716 15202 30772 15214
rect 30716 15150 30718 15202
rect 30770 15150 30772 15202
rect 30716 15148 30772 15150
rect 31164 15148 31220 15262
rect 30716 15092 31220 15148
rect 31276 15316 31332 15326
rect 31052 14420 31108 15092
rect 31276 14530 31332 15260
rect 31276 14478 31278 14530
rect 31330 14478 31332 14530
rect 31052 14364 31220 14420
rect 30604 14028 30996 14084
rect 29484 12798 29486 12850
rect 29538 12798 29540 12850
rect 29484 12786 29540 12798
rect 29708 13356 30100 13412
rect 30268 13746 30324 13758
rect 30268 13694 30270 13746
rect 30322 13694 30324 13746
rect 29708 12516 29764 13356
rect 29596 12460 29764 12516
rect 30044 12852 30100 12862
rect 30268 12852 30324 13694
rect 30044 12850 30324 12852
rect 30044 12798 30046 12850
rect 30098 12798 30324 12850
rect 30044 12796 30324 12798
rect 29260 12236 29428 12292
rect 29260 12068 29316 12078
rect 29260 11974 29316 12012
rect 29372 11620 29428 12236
rect 29260 11564 29428 11620
rect 29596 12290 29652 12460
rect 29596 12238 29598 12290
rect 29650 12238 29652 12290
rect 29260 11284 29316 11564
rect 29596 11508 29652 12238
rect 29596 11442 29652 11452
rect 29708 12290 29764 12302
rect 29708 12238 29710 12290
rect 29762 12238 29764 12290
rect 29708 12068 29764 12238
rect 30044 12292 30100 12796
rect 30380 12738 30436 14028
rect 30492 14018 30548 14028
rect 30492 13860 30548 13870
rect 30492 13766 30548 13804
rect 30604 13748 30660 13758
rect 30604 13654 30660 13692
rect 30828 13186 30884 13198
rect 30828 13134 30830 13186
rect 30882 13134 30884 13186
rect 30828 12740 30884 13134
rect 30380 12686 30382 12738
rect 30434 12686 30436 12738
rect 30380 12674 30436 12686
rect 30716 12684 30884 12740
rect 30044 12226 30100 12236
rect 30268 12292 30324 12302
rect 30268 12198 30324 12236
rect 29932 12180 29988 12190
rect 29932 12086 29988 12124
rect 30492 12180 30548 12190
rect 30492 12086 30548 12124
rect 29260 10834 29316 11228
rect 29260 10782 29262 10834
rect 29314 10782 29316 10834
rect 29260 10770 29316 10782
rect 29372 11394 29428 11406
rect 29372 11342 29374 11394
rect 29426 11342 29428 11394
rect 29148 10434 29204 10444
rect 28924 10332 29092 10388
rect 28812 9268 28868 9278
rect 28252 9266 28532 9268
rect 28252 9214 28254 9266
rect 28306 9214 28532 9266
rect 28252 9212 28532 9214
rect 28700 9266 28868 9268
rect 28700 9214 28814 9266
rect 28866 9214 28868 9266
rect 28700 9212 28868 9214
rect 28252 9202 28308 9212
rect 26908 8258 27412 8260
rect 26908 8206 26910 8258
rect 26962 8206 27412 8258
rect 26908 8204 27412 8206
rect 26460 6692 26516 6702
rect 26236 6514 26292 6524
rect 26348 6578 26404 6590
rect 26348 6526 26350 6578
rect 26402 6526 26404 6578
rect 26348 6356 26404 6526
rect 26460 6466 26516 6636
rect 26684 6580 26740 6860
rect 26460 6414 26462 6466
rect 26514 6414 26516 6466
rect 26460 6402 26516 6414
rect 26572 6524 26740 6580
rect 26796 6690 26852 6702
rect 26796 6638 26798 6690
rect 26850 6638 26852 6690
rect 26348 6290 26404 6300
rect 26236 6244 26292 6254
rect 26236 5908 26292 6188
rect 26348 5908 26404 5918
rect 26236 5906 26404 5908
rect 26236 5854 26350 5906
rect 26402 5854 26404 5906
rect 26236 5852 26404 5854
rect 25900 5814 25956 5852
rect 26348 5842 26404 5852
rect 25788 5516 25956 5572
rect 25788 5348 25844 5358
rect 25676 5236 25732 5246
rect 25788 5236 25844 5292
rect 25676 5234 25844 5236
rect 25676 5182 25678 5234
rect 25730 5182 25844 5234
rect 25676 5180 25844 5182
rect 25676 5170 25732 5180
rect 25900 5122 25956 5516
rect 25900 5070 25902 5122
rect 25954 5070 25956 5122
rect 25900 5058 25956 5070
rect 26012 5180 26404 5236
rect 26012 5122 26068 5180
rect 26012 5070 26014 5122
rect 26066 5070 26068 5122
rect 25564 4386 25620 4396
rect 25564 4228 25620 4238
rect 26012 4228 26068 5070
rect 26348 5122 26404 5180
rect 26348 5070 26350 5122
rect 26402 5070 26404 5122
rect 26348 5058 26404 5070
rect 26572 5012 26628 6524
rect 26796 6468 26852 6638
rect 26684 6412 26796 6468
rect 26684 6130 26740 6412
rect 26796 6402 26852 6412
rect 26684 6078 26686 6130
rect 26738 6078 26740 6130
rect 26684 6020 26740 6078
rect 26684 5954 26740 5964
rect 26908 6130 26964 8204
rect 27244 8036 27300 8046
rect 27244 7942 27300 7980
rect 27356 7698 27412 8204
rect 27356 7646 27358 7698
rect 27410 7646 27412 7698
rect 27356 7634 27412 7646
rect 27580 8148 27636 8158
rect 27580 7476 27636 8092
rect 27804 8146 27860 8876
rect 27916 8372 27972 8382
rect 28252 8372 28308 8382
rect 27916 8370 28308 8372
rect 27916 8318 27918 8370
rect 27970 8318 28254 8370
rect 28306 8318 28308 8370
rect 27916 8316 28308 8318
rect 27916 8306 27972 8316
rect 28252 8306 28308 8316
rect 27804 8094 27806 8146
rect 27858 8094 27860 8146
rect 27804 7700 27860 8094
rect 28364 8148 28420 8158
rect 28364 8054 28420 8092
rect 28476 8146 28532 9212
rect 28812 8818 28868 9212
rect 28812 8766 28814 8818
rect 28866 8766 28868 8818
rect 28812 8754 28868 8766
rect 28476 8094 28478 8146
rect 28530 8094 28532 8146
rect 28476 8036 28532 8094
rect 28476 7970 28532 7980
rect 28252 7700 28308 7710
rect 28924 7700 28980 10332
rect 29148 9828 29204 9838
rect 29148 9734 29204 9772
rect 29372 9268 29428 11342
rect 29596 9940 29652 9950
rect 29708 9940 29764 12012
rect 30716 11956 30772 12684
rect 30828 12404 30884 12414
rect 30940 12404 30996 14028
rect 31052 13860 31108 13870
rect 31052 13766 31108 13804
rect 31052 12740 31108 12750
rect 31164 12740 31220 14364
rect 31276 14084 31332 14478
rect 31276 14018 31332 14028
rect 31388 13860 31444 16044
rect 31500 14868 31556 17500
rect 31724 17462 31780 17500
rect 31836 16882 31892 16894
rect 31836 16830 31838 16882
rect 31890 16830 31892 16882
rect 31836 16660 31892 16830
rect 31836 16594 31892 16604
rect 31612 15874 31668 15886
rect 31612 15822 31614 15874
rect 31666 15822 31668 15874
rect 31612 15652 31668 15822
rect 31612 15586 31668 15596
rect 31724 15876 31780 15886
rect 31724 15426 31780 15820
rect 31724 15374 31726 15426
rect 31778 15374 31780 15426
rect 31500 14802 31556 14812
rect 31612 15314 31668 15326
rect 31612 15262 31614 15314
rect 31666 15262 31668 15314
rect 31108 12684 31220 12740
rect 31276 13804 31444 13860
rect 31500 14642 31556 14654
rect 31500 14590 31502 14642
rect 31554 14590 31556 14642
rect 31052 12516 31108 12684
rect 31052 12450 31108 12460
rect 30828 12402 30940 12404
rect 30828 12350 30830 12402
rect 30882 12350 30940 12402
rect 30828 12348 30940 12350
rect 30828 12338 30884 12348
rect 30940 12310 30996 12348
rect 31052 12292 31108 12302
rect 31276 12292 31332 13804
rect 31388 13634 31444 13646
rect 31388 13582 31390 13634
rect 31442 13582 31444 13634
rect 31388 12740 31444 13582
rect 31500 12964 31556 14590
rect 31612 13522 31668 15262
rect 31724 14418 31780 15374
rect 31724 14366 31726 14418
rect 31778 14366 31780 14418
rect 31724 14354 31780 14366
rect 31836 14868 31892 14878
rect 31612 13470 31614 13522
rect 31666 13470 31668 13522
rect 31612 13186 31668 13470
rect 31612 13134 31614 13186
rect 31666 13134 31668 13186
rect 31612 13122 31668 13134
rect 31500 12908 31668 12964
rect 31388 12674 31444 12684
rect 31500 12738 31556 12750
rect 31500 12686 31502 12738
rect 31554 12686 31556 12738
rect 31500 12628 31556 12686
rect 31500 12562 31556 12572
rect 31052 12290 31332 12292
rect 31052 12238 31054 12290
rect 31106 12238 31332 12290
rect 31052 12236 31332 12238
rect 31388 12404 31444 12414
rect 31388 12292 31444 12348
rect 31500 12292 31556 12302
rect 31388 12290 31556 12292
rect 31388 12238 31502 12290
rect 31554 12238 31556 12290
rect 31388 12236 31556 12238
rect 31052 12180 31108 12236
rect 31500 12226 31556 12236
rect 31052 12114 31108 12124
rect 30492 11900 30772 11956
rect 31164 11956 31220 11966
rect 30156 11732 30212 11742
rect 30156 11620 30212 11676
rect 30156 11564 30324 11620
rect 30156 11394 30212 11406
rect 30156 11342 30158 11394
rect 30210 11342 30212 11394
rect 29932 11284 29988 11294
rect 29596 9938 29764 9940
rect 29596 9886 29598 9938
rect 29650 9886 29764 9938
rect 29596 9884 29764 9886
rect 29820 11228 29932 11284
rect 29596 9492 29652 9884
rect 29820 9716 29876 11228
rect 29932 11218 29988 11228
rect 30156 11060 30212 11342
rect 30268 11282 30324 11564
rect 30268 11230 30270 11282
rect 30322 11230 30324 11282
rect 30268 11218 30324 11230
rect 29932 11004 30212 11060
rect 29932 10610 29988 11004
rect 30156 10836 30212 10846
rect 30156 10742 30212 10780
rect 29932 10558 29934 10610
rect 29986 10558 29988 10610
rect 29932 10388 29988 10558
rect 30044 10500 30100 10510
rect 30044 10406 30100 10444
rect 29932 10322 29988 10332
rect 30268 10052 30324 10062
rect 29820 9660 29988 9716
rect 29596 9426 29652 9436
rect 29372 9202 29428 9212
rect 29260 9156 29316 9166
rect 29260 9062 29316 9100
rect 29708 9156 29764 9166
rect 29484 8818 29540 8830
rect 29484 8766 29486 8818
rect 29538 8766 29540 8818
rect 27804 7698 28252 7700
rect 27804 7646 27806 7698
rect 27858 7646 28252 7698
rect 27804 7644 28252 7646
rect 27804 7634 27860 7644
rect 28252 7606 28308 7644
rect 28812 7644 28980 7700
rect 29036 8258 29092 8270
rect 29036 8206 29038 8258
rect 29090 8206 29092 8258
rect 29036 7700 29092 8206
rect 29484 8258 29540 8766
rect 29484 8206 29486 8258
rect 29538 8206 29540 8258
rect 29484 8194 29540 8206
rect 29708 8146 29764 9100
rect 29708 8094 29710 8146
rect 29762 8094 29764 8146
rect 29708 8082 29764 8094
rect 29596 8036 29652 8046
rect 29596 7942 29652 7980
rect 27580 7410 27636 7420
rect 28028 7364 28084 7374
rect 26908 6078 26910 6130
rect 26962 6078 26964 6130
rect 26908 6020 26964 6078
rect 26908 5954 26964 5964
rect 27244 7028 27300 7038
rect 27132 5908 27188 5918
rect 27020 5906 27188 5908
rect 27020 5854 27134 5906
rect 27186 5854 27188 5906
rect 27020 5852 27188 5854
rect 27020 5794 27076 5852
rect 27132 5842 27188 5852
rect 27020 5742 27022 5794
rect 27074 5742 27076 5794
rect 27020 5730 27076 5742
rect 27244 5684 27300 6972
rect 27468 6690 27524 6702
rect 27468 6638 27470 6690
rect 27522 6638 27524 6690
rect 27468 6132 27524 6638
rect 27468 6066 27524 6076
rect 27132 5628 27300 5684
rect 27692 6020 27748 6030
rect 26908 5572 26964 5582
rect 26908 5234 26964 5516
rect 26908 5182 26910 5234
rect 26962 5182 26964 5234
rect 26908 5170 26964 5182
rect 27020 5236 27076 5246
rect 27020 5122 27076 5180
rect 27020 5070 27022 5122
rect 27074 5070 27076 5122
rect 27020 5058 27076 5070
rect 26796 5012 26852 5022
rect 26460 5010 26852 5012
rect 26460 4958 26798 5010
rect 26850 4958 26852 5010
rect 26460 4956 26852 4958
rect 26460 4676 26516 4956
rect 26796 4946 26852 4956
rect 26236 4620 26516 4676
rect 26236 4562 26292 4620
rect 26236 4510 26238 4562
rect 26290 4510 26292 4562
rect 26236 4498 26292 4510
rect 25564 4226 26068 4228
rect 25564 4174 25566 4226
rect 25618 4174 26068 4226
rect 25564 4172 26068 4174
rect 25564 4162 25620 4172
rect 25004 2818 25060 2828
rect 16604 2594 16660 2604
rect 27132 2660 27188 5628
rect 27692 5236 27748 5964
rect 28028 6018 28084 7308
rect 28812 7362 28868 7644
rect 29036 7634 29092 7644
rect 28812 7310 28814 7362
rect 28866 7310 28868 7362
rect 28364 6802 28420 6814
rect 28364 6750 28366 6802
rect 28418 6750 28420 6802
rect 28028 5966 28030 6018
rect 28082 5966 28084 6018
rect 28028 5954 28084 5966
rect 28140 6580 28196 6590
rect 28140 5908 28196 6524
rect 28364 6580 28420 6750
rect 28812 6804 28868 7310
rect 28476 6692 28532 6702
rect 28476 6598 28532 6636
rect 28364 6514 28420 6524
rect 28812 6468 28868 6748
rect 28812 6402 28868 6412
rect 28924 7474 28980 7486
rect 28924 7422 28926 7474
rect 28978 7422 28980 7474
rect 28140 5814 28196 5852
rect 27804 5794 27860 5806
rect 27804 5742 27806 5794
rect 27858 5742 27860 5794
rect 27804 5348 27860 5742
rect 28924 5684 28980 7422
rect 29708 7476 29764 7486
rect 29260 6804 29316 6814
rect 29260 6710 29316 6748
rect 29036 6020 29092 6030
rect 29708 6020 29764 7420
rect 29820 7250 29876 7262
rect 29820 7198 29822 7250
rect 29874 7198 29876 7250
rect 29820 6804 29876 7198
rect 29820 6738 29876 6748
rect 29932 6132 29988 9660
rect 30268 8484 30324 9996
rect 30268 8418 30324 8428
rect 30044 8148 30100 8158
rect 30044 7474 30100 8092
rect 30380 8148 30436 8158
rect 30380 8054 30436 8092
rect 30156 8036 30212 8046
rect 30156 7942 30212 7980
rect 30044 7422 30046 7474
rect 30098 7422 30100 7474
rect 30044 7410 30100 7422
rect 29932 6038 29988 6076
rect 29820 6020 29876 6030
rect 29708 6018 29876 6020
rect 29708 5966 29822 6018
rect 29874 5966 29876 6018
rect 29708 5964 29876 5966
rect 29036 5906 29092 5964
rect 29820 5954 29876 5964
rect 29036 5854 29038 5906
rect 29090 5854 29092 5906
rect 29036 5842 29092 5854
rect 29372 5908 29428 5918
rect 29372 5794 29428 5852
rect 29372 5742 29374 5794
rect 29426 5742 29428 5794
rect 29372 5730 29428 5742
rect 29932 5684 29988 5694
rect 28812 5628 28980 5684
rect 29596 5682 29988 5684
rect 29596 5630 29934 5682
rect 29986 5630 29988 5682
rect 29596 5628 29988 5630
rect 27804 5282 27860 5292
rect 28476 5460 28532 5470
rect 27244 5234 27748 5236
rect 27244 5182 27694 5234
rect 27746 5182 27748 5234
rect 27244 5180 27748 5182
rect 27244 4562 27300 5180
rect 27692 5170 27748 5180
rect 28140 5234 28196 5246
rect 28140 5182 28142 5234
rect 28194 5182 28196 5234
rect 28140 5012 28196 5182
rect 28476 5124 28532 5404
rect 28476 5030 28532 5068
rect 28812 5348 28868 5628
rect 29596 5460 29652 5628
rect 29932 5618 29988 5628
rect 28140 4788 28196 4956
rect 28140 4722 28196 4732
rect 27244 4510 27246 4562
rect 27298 4510 27300 4562
rect 27244 4498 27300 4510
rect 28812 4562 28868 5292
rect 28812 4510 28814 4562
rect 28866 4510 28868 4562
rect 28812 4498 28868 4510
rect 28924 5404 29652 5460
rect 28924 4450 28980 5404
rect 29148 5236 29204 5246
rect 29148 5122 29204 5180
rect 30380 5236 30436 5246
rect 30380 5142 30436 5180
rect 29148 5070 29150 5122
rect 29202 5070 29204 5122
rect 29148 5058 29204 5070
rect 29484 5124 29540 5134
rect 29372 5010 29428 5022
rect 29372 4958 29374 5010
rect 29426 4958 29428 5010
rect 29372 4676 29428 4958
rect 28924 4398 28926 4450
rect 28978 4398 28980 4450
rect 28924 4386 28980 4398
rect 29036 4620 29428 4676
rect 28812 4116 28868 4126
rect 29036 4116 29092 4620
rect 29484 4562 29540 5068
rect 29708 5012 29764 5022
rect 29708 4918 29764 4956
rect 29484 4510 29486 4562
rect 29538 4510 29540 4562
rect 29484 4498 29540 4510
rect 30380 4564 30436 4574
rect 30380 4470 30436 4508
rect 28812 4114 29092 4116
rect 28812 4062 28814 4114
rect 28866 4062 29092 4114
rect 28812 4060 29092 4062
rect 28812 4050 28868 4060
rect 28812 3668 28868 3678
rect 28868 3612 29092 3668
rect 28812 3574 28868 3612
rect 29036 3554 29092 3612
rect 29036 3502 29038 3554
rect 29090 3502 29092 3554
rect 29036 3490 29092 3502
rect 27132 2594 27188 2604
rect 28924 3444 28980 3454
rect 28924 800 28980 3388
rect 30044 3444 30100 3454
rect 30044 3330 30100 3388
rect 30044 3278 30046 3330
rect 30098 3278 30100 3330
rect 30044 3266 30100 3278
rect 30492 1652 30548 11900
rect 31164 11862 31220 11900
rect 31388 11508 31444 11518
rect 31388 11414 31444 11452
rect 31052 11396 31108 11406
rect 31052 11302 31108 11340
rect 30940 11284 30996 11294
rect 30940 11190 30996 11228
rect 30604 10724 30660 10734
rect 30604 10610 30660 10668
rect 30604 10558 30606 10610
rect 30658 10558 30660 10610
rect 30604 10546 30660 10558
rect 31500 10722 31556 10734
rect 31500 10670 31502 10722
rect 31554 10670 31556 10722
rect 31276 10500 31332 10510
rect 31276 10406 31332 10444
rect 30940 10388 30996 10398
rect 30828 10386 30996 10388
rect 30828 10334 30942 10386
rect 30994 10334 30996 10386
rect 30828 10332 30996 10334
rect 30604 6132 30660 6142
rect 30604 6038 30660 6076
rect 30716 4676 30772 4686
rect 30716 4562 30772 4620
rect 30716 4510 30718 4562
rect 30770 4510 30772 4562
rect 30716 4498 30772 4510
rect 30828 4562 30884 10332
rect 30940 10322 30996 10332
rect 31500 9268 31556 10670
rect 31612 9828 31668 12908
rect 31836 10948 31892 14812
rect 32172 14532 32228 17614
rect 32732 17666 32788 18172
rect 32732 17614 32734 17666
rect 32786 17614 32788 17666
rect 32732 17108 32788 17614
rect 32508 17052 32788 17108
rect 32508 16994 32564 17052
rect 32508 16942 32510 16994
rect 32562 16942 32564 16994
rect 32508 16930 32564 16942
rect 32956 15988 33012 22876
rect 33068 22866 33124 22876
rect 33404 22482 33460 22494
rect 33404 22430 33406 22482
rect 33458 22430 33460 22482
rect 33068 21586 33124 21598
rect 33068 21534 33070 21586
rect 33122 21534 33124 21586
rect 33068 20018 33124 21534
rect 33292 21586 33348 21598
rect 33292 21534 33294 21586
rect 33346 21534 33348 21586
rect 33292 20244 33348 21534
rect 33292 20130 33348 20188
rect 33292 20078 33294 20130
rect 33346 20078 33348 20130
rect 33292 20066 33348 20078
rect 33068 19966 33070 20018
rect 33122 19966 33124 20018
rect 33068 19348 33124 19966
rect 33068 19282 33124 19292
rect 33404 18004 33460 22430
rect 33516 22484 33572 22988
rect 33516 22418 33572 22428
rect 33852 22370 33908 24668
rect 33852 22318 33854 22370
rect 33906 22318 33908 22370
rect 33852 22306 33908 22318
rect 33964 24612 34020 25228
rect 34076 25218 34132 25228
rect 33852 21924 33908 21934
rect 33852 21810 33908 21868
rect 33852 21758 33854 21810
rect 33906 21758 33908 21810
rect 33852 21746 33908 21758
rect 33516 21586 33572 21598
rect 33516 21534 33518 21586
rect 33570 21534 33572 21586
rect 33516 21252 33572 21534
rect 33516 20802 33572 21196
rect 33516 20750 33518 20802
rect 33570 20750 33572 20802
rect 33516 20468 33572 20750
rect 33516 20402 33572 20412
rect 33740 21586 33796 21598
rect 33740 21534 33742 21586
rect 33794 21534 33796 21586
rect 33628 20132 33684 20142
rect 33628 19796 33684 20076
rect 33628 19730 33684 19740
rect 33740 19684 33796 21534
rect 33852 21588 33908 21598
rect 33852 21026 33908 21532
rect 33852 20974 33854 21026
rect 33906 20974 33908 21026
rect 33852 20580 33908 20974
rect 33852 20514 33908 20524
rect 33964 20188 34020 24556
rect 34412 23828 34468 25454
rect 35084 25506 35140 25518
rect 35084 25454 35086 25506
rect 35138 25454 35140 25506
rect 34972 24722 35028 24734
rect 34972 24670 34974 24722
rect 35026 24670 35028 24722
rect 34972 24612 35028 24670
rect 34972 24546 35028 24556
rect 34524 23828 34580 23838
rect 34412 23826 34580 23828
rect 34412 23774 34526 23826
rect 34578 23774 34580 23826
rect 34412 23772 34580 23774
rect 34524 23762 34580 23772
rect 35084 23714 35140 25454
rect 35532 25506 35588 25518
rect 35532 25454 35534 25506
rect 35586 25454 35588 25506
rect 35532 24722 35588 25454
rect 35532 24670 35534 24722
rect 35586 24670 35588 24722
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35532 23940 35588 24670
rect 35084 23662 35086 23714
rect 35138 23662 35140 23714
rect 34860 23156 34916 23166
rect 34300 23044 34356 23054
rect 34300 22950 34356 22988
rect 34860 23042 34916 23100
rect 35084 23154 35140 23662
rect 35084 23102 35086 23154
rect 35138 23102 35140 23154
rect 35084 23090 35140 23102
rect 35196 23884 35588 23940
rect 35756 25394 35812 25406
rect 35756 25342 35758 25394
rect 35810 25342 35812 25394
rect 35196 23156 35252 23884
rect 35756 23716 35812 25342
rect 36204 25284 36260 25294
rect 36204 25190 36260 25228
rect 36988 25284 37044 25294
rect 36988 25190 37044 25228
rect 36092 24834 36148 24846
rect 36092 24782 36094 24834
rect 36146 24782 36148 24834
rect 35756 23650 35812 23660
rect 35980 24610 36036 24622
rect 35980 24558 35982 24610
rect 36034 24558 36036 24610
rect 35196 23090 35252 23100
rect 35756 23154 35812 23166
rect 35756 23102 35758 23154
rect 35810 23102 35812 23154
rect 34860 22990 34862 23042
rect 34914 22990 34916 23042
rect 34860 22978 34916 22990
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35196 22482 35252 22494
rect 35196 22430 35198 22482
rect 35250 22430 35252 22482
rect 34524 22372 34580 22382
rect 33628 19012 33684 19022
rect 33740 19012 33796 19628
rect 33628 19010 33796 19012
rect 33628 18958 33630 19010
rect 33682 18958 33796 19010
rect 33628 18956 33796 18958
rect 33628 18946 33684 18956
rect 33404 17938 33460 17948
rect 33404 17556 33460 17566
rect 33404 17462 33460 17500
rect 33740 16884 33796 18956
rect 33852 20132 34020 20188
rect 34076 21586 34132 21598
rect 34076 21534 34078 21586
rect 34130 21534 34132 21586
rect 34076 20132 34132 21534
rect 34524 20356 34580 22316
rect 34972 22370 35028 22382
rect 34972 22318 34974 22370
rect 35026 22318 35028 22370
rect 34972 21812 35028 22318
rect 34972 21746 35028 21756
rect 35196 21810 35252 22430
rect 35756 22370 35812 23102
rect 35980 23156 36036 24558
rect 36092 23940 36148 24782
rect 36876 24722 36932 24734
rect 36876 24670 36878 24722
rect 36930 24670 36932 24722
rect 36876 24612 36932 24670
rect 36876 24546 36932 24556
rect 36092 23874 36148 23884
rect 35980 23090 36036 23100
rect 36988 23716 37044 23726
rect 36204 22484 36260 22522
rect 36204 22418 36260 22428
rect 35756 22318 35758 22370
rect 35810 22318 35812 22370
rect 35756 22306 35812 22318
rect 35980 22372 36036 22382
rect 35980 22278 36036 22316
rect 35196 21758 35198 21810
rect 35250 21758 35252 21810
rect 35196 21746 35252 21758
rect 36204 22260 36260 22270
rect 35084 21698 35140 21710
rect 35084 21646 35086 21698
rect 35138 21646 35140 21698
rect 34972 21588 35028 21598
rect 34748 21586 35028 21588
rect 34748 21534 34974 21586
rect 35026 21534 35028 21586
rect 34748 21532 35028 21534
rect 34636 21476 34692 21486
rect 34636 21382 34692 21420
rect 34748 20916 34804 21532
rect 34972 21522 35028 21532
rect 35084 21588 35140 21646
rect 35084 21522 35140 21532
rect 35644 21588 35700 21598
rect 35084 21364 35140 21374
rect 35084 20916 35140 21308
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35644 21026 35700 21532
rect 35644 20974 35646 21026
rect 35698 20974 35700 21026
rect 35644 20962 35700 20974
rect 34636 20804 34692 20814
rect 34748 20804 34804 20860
rect 34636 20802 34804 20804
rect 34636 20750 34638 20802
rect 34690 20750 34804 20802
rect 34636 20748 34804 20750
rect 34636 20738 34692 20748
rect 34748 20356 34804 20748
rect 34524 20300 34692 20356
rect 33852 17108 33908 20132
rect 34076 20066 34132 20076
rect 34524 20130 34580 20142
rect 34524 20078 34526 20130
rect 34578 20078 34580 20130
rect 34524 20020 34580 20078
rect 34300 19908 34356 19918
rect 34300 19814 34356 19852
rect 33964 19012 34020 19022
rect 33964 18918 34020 18956
rect 34524 19012 34580 19964
rect 34524 18946 34580 18956
rect 34636 18116 34692 20300
rect 34748 20290 34804 20300
rect 34860 20860 35140 20916
rect 34860 20242 34916 20860
rect 35084 20802 35140 20860
rect 35868 20916 35924 20926
rect 35868 20822 35924 20860
rect 36204 20914 36260 22204
rect 36988 22146 37044 23660
rect 36988 22094 36990 22146
rect 37042 22094 37044 22146
rect 36988 22082 37044 22094
rect 36204 20862 36206 20914
rect 36258 20862 36260 20914
rect 36204 20850 36260 20862
rect 36316 21588 36372 21598
rect 35084 20750 35086 20802
rect 35138 20750 35140 20802
rect 35084 20738 35140 20750
rect 36316 20802 36372 21532
rect 36316 20750 36318 20802
rect 36370 20750 36372 20802
rect 36316 20738 36372 20750
rect 34860 20190 34862 20242
rect 34914 20190 34916 20242
rect 34860 20178 34916 20190
rect 34972 20690 35028 20702
rect 34972 20638 34974 20690
rect 35026 20638 35028 20690
rect 34972 20132 35028 20638
rect 36092 20578 36148 20590
rect 36092 20526 36094 20578
rect 36146 20526 36148 20578
rect 36092 20188 36148 20526
rect 36092 20132 36708 20188
rect 34972 20066 35028 20076
rect 36204 20130 36260 20132
rect 36204 20078 36206 20130
rect 36258 20078 36260 20130
rect 36204 20066 36260 20078
rect 35980 20018 36036 20030
rect 35980 19966 35982 20018
rect 36034 19966 36036 20018
rect 35980 19796 36036 19966
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35868 19010 35924 19022
rect 35868 18958 35870 19010
rect 35922 18958 35924 19010
rect 35868 18564 35924 18958
rect 35644 18508 35924 18564
rect 35532 18452 35588 18462
rect 35644 18452 35700 18508
rect 35532 18450 35700 18452
rect 35532 18398 35534 18450
rect 35586 18398 35700 18450
rect 35532 18396 35700 18398
rect 34636 18060 34916 18116
rect 34300 18004 34356 18014
rect 34356 17948 34468 18004
rect 34300 17938 34356 17948
rect 34300 17668 34356 17678
rect 34300 17574 34356 17612
rect 34076 17556 34132 17566
rect 33852 17052 34020 17108
rect 33852 16884 33908 16894
rect 33740 16882 33908 16884
rect 33740 16830 33854 16882
rect 33906 16830 33908 16882
rect 33740 16828 33908 16830
rect 33404 16212 33460 16222
rect 33404 16100 33460 16156
rect 32956 15922 33012 15932
rect 33068 16098 33460 16100
rect 33068 16046 33406 16098
rect 33458 16046 33460 16098
rect 33068 16044 33460 16046
rect 32956 15316 33012 15326
rect 32956 15222 33012 15260
rect 32172 14466 32228 14476
rect 32396 14644 32452 14654
rect 31948 14420 32004 14430
rect 31948 13972 32004 14364
rect 31948 13970 32228 13972
rect 31948 13918 31950 13970
rect 32002 13918 32228 13970
rect 31948 13916 32228 13918
rect 31948 13906 32004 13916
rect 32172 12962 32228 13916
rect 32172 12910 32174 12962
rect 32226 12910 32228 12962
rect 32172 12898 32228 12910
rect 32284 13748 32340 13758
rect 31724 10892 31892 10948
rect 31724 10052 31780 10892
rect 31836 10724 31892 10734
rect 31836 10630 31892 10668
rect 31724 9986 31780 9996
rect 31612 9772 31780 9828
rect 31500 9202 31556 9212
rect 31612 9604 31668 9614
rect 31612 9042 31668 9548
rect 31612 8990 31614 9042
rect 31666 8990 31668 9042
rect 31612 8978 31668 8990
rect 31724 8260 31780 9772
rect 31388 8204 31724 8260
rect 31388 6690 31444 8204
rect 31724 8194 31780 8204
rect 31948 9042 32004 9054
rect 31948 8990 31950 9042
rect 32002 8990 32004 9042
rect 31948 8036 32004 8990
rect 32060 8260 32116 8298
rect 32060 8194 32116 8204
rect 32172 8148 32228 8158
rect 32284 8148 32340 13692
rect 32396 13074 32452 14588
rect 33068 13860 33124 16044
rect 33404 16034 33460 16044
rect 33516 16100 33572 16110
rect 33516 16006 33572 16044
rect 33628 15988 33684 15998
rect 33180 15876 33236 15886
rect 33180 15782 33236 15820
rect 33628 15652 33684 15932
rect 33180 15596 33684 15652
rect 33180 14530 33236 15596
rect 33404 15314 33460 15326
rect 33404 15262 33406 15314
rect 33458 15262 33460 15314
rect 33404 15204 33460 15262
rect 33628 15314 33684 15326
rect 33628 15262 33630 15314
rect 33682 15262 33684 15314
rect 33404 15138 33460 15148
rect 33516 15202 33572 15214
rect 33516 15150 33518 15202
rect 33570 15150 33572 15202
rect 33180 14478 33182 14530
rect 33234 14478 33236 14530
rect 33180 14466 33236 14478
rect 33404 14980 33460 14990
rect 33292 14196 33348 14206
rect 33292 13970 33348 14140
rect 33292 13918 33294 13970
rect 33346 13918 33348 13970
rect 33292 13906 33348 13918
rect 33180 13860 33236 13870
rect 33068 13858 33236 13860
rect 33068 13806 33182 13858
rect 33234 13806 33236 13858
rect 33068 13804 33236 13806
rect 33180 13794 33236 13804
rect 32508 13636 32564 13646
rect 32508 13186 32564 13580
rect 32508 13134 32510 13186
rect 32562 13134 32564 13186
rect 32508 13122 32564 13134
rect 32396 13022 32398 13074
rect 32450 13022 32452 13074
rect 32396 13010 32452 13022
rect 33292 12404 33348 12414
rect 33404 12404 33460 14924
rect 33516 14756 33572 15150
rect 33516 14690 33572 14700
rect 33628 14644 33684 15262
rect 33740 14980 33796 16828
rect 33852 16818 33908 16828
rect 33964 16212 34020 17052
rect 33964 16146 34020 16156
rect 34076 16882 34132 17500
rect 34412 17108 34468 17948
rect 34524 17890 34580 17902
rect 34524 17838 34526 17890
rect 34578 17838 34580 17890
rect 34524 17556 34580 17838
rect 34748 17892 34804 17902
rect 34748 17778 34804 17836
rect 34748 17726 34750 17778
rect 34802 17726 34804 17778
rect 34748 17714 34804 17726
rect 34524 17490 34580 17500
rect 34412 17052 34580 17108
rect 34076 16830 34078 16882
rect 34130 16830 34132 16882
rect 34076 15988 34132 16830
rect 34412 16884 34468 16894
rect 34412 16790 34468 16828
rect 34412 16212 34468 16222
rect 34300 16100 34356 16110
rect 34300 16006 34356 16044
rect 34076 15922 34132 15932
rect 34076 15540 34132 15550
rect 33740 14914 33796 14924
rect 33964 15204 34020 15214
rect 33852 14756 33908 14766
rect 33628 14578 33684 14588
rect 33740 14754 33908 14756
rect 33740 14702 33854 14754
rect 33906 14702 33908 14754
rect 33740 14700 33908 14702
rect 33628 14420 33684 14430
rect 33628 14326 33684 14364
rect 33628 13860 33684 13870
rect 33740 13860 33796 14700
rect 33852 14690 33908 14700
rect 33684 13804 33796 13860
rect 33628 13766 33684 13804
rect 33852 13748 33908 13758
rect 33852 13654 33908 13692
rect 33292 12402 33460 12404
rect 33292 12350 33294 12402
rect 33346 12350 33460 12402
rect 33292 12348 33460 12350
rect 33292 12338 33348 12348
rect 33180 12178 33236 12190
rect 33180 12126 33182 12178
rect 33234 12126 33236 12178
rect 32956 11620 33012 11630
rect 33180 11620 33236 12126
rect 33852 12068 33908 12078
rect 33740 12066 33908 12068
rect 33740 12014 33854 12066
rect 33906 12014 33908 12066
rect 33740 12012 33908 12014
rect 33012 11564 33236 11620
rect 33292 11954 33348 11966
rect 33292 11902 33294 11954
rect 33346 11902 33348 11954
rect 32956 11170 33012 11564
rect 33292 11394 33348 11902
rect 33740 11620 33796 12012
rect 33852 12002 33908 12012
rect 33740 11506 33796 11564
rect 33740 11454 33742 11506
rect 33794 11454 33796 11506
rect 33740 11442 33796 11454
rect 33292 11342 33294 11394
rect 33346 11342 33348 11394
rect 33292 11330 33348 11342
rect 33516 11396 33572 11406
rect 32956 11118 32958 11170
rect 33010 11118 33012 11170
rect 32956 10276 33012 11118
rect 33516 10610 33572 11340
rect 33740 10948 33796 10958
rect 33516 10558 33518 10610
rect 33570 10558 33572 10610
rect 33516 10546 33572 10558
rect 33628 10724 33684 10734
rect 33180 10388 33236 10398
rect 33180 10386 33460 10388
rect 33180 10334 33182 10386
rect 33234 10334 33460 10386
rect 33180 10332 33460 10334
rect 33180 10322 33236 10332
rect 32956 10210 33012 10220
rect 32620 10052 32676 10062
rect 32396 9602 32452 9614
rect 32396 9550 32398 9602
rect 32450 9550 32452 9602
rect 32396 9268 32452 9550
rect 32396 9202 32452 9212
rect 32508 8932 32564 8942
rect 32508 8838 32564 8876
rect 32172 8146 32340 8148
rect 32172 8094 32174 8146
rect 32226 8094 32340 8146
rect 32172 8092 32340 8094
rect 32060 8036 32116 8046
rect 31948 7980 32060 8036
rect 31948 7588 32004 7598
rect 31948 7362 32004 7532
rect 32060 7474 32116 7980
rect 32060 7422 32062 7474
rect 32114 7422 32116 7474
rect 32060 7410 32116 7422
rect 31948 7310 31950 7362
rect 32002 7310 32004 7362
rect 31948 7298 32004 7310
rect 31388 6638 31390 6690
rect 31442 6638 31444 6690
rect 31388 6626 31444 6638
rect 31612 6692 31668 6702
rect 31612 6598 31668 6636
rect 32060 6692 32116 6702
rect 32172 6692 32228 8092
rect 32508 7588 32564 7598
rect 32508 7494 32564 7532
rect 32620 7028 32676 9996
rect 33404 9826 33460 10332
rect 33404 9774 33406 9826
rect 33458 9774 33460 9826
rect 33404 9762 33460 9774
rect 33516 9602 33572 9614
rect 33516 9550 33518 9602
rect 33570 9550 33572 9602
rect 33516 9380 33572 9550
rect 33628 9602 33684 10668
rect 33740 10722 33796 10892
rect 33740 10670 33742 10722
rect 33794 10670 33796 10722
rect 33740 10658 33796 10670
rect 33628 9550 33630 9602
rect 33682 9550 33684 9602
rect 33628 9538 33684 9550
rect 33516 9324 33684 9380
rect 32732 8146 32788 8158
rect 32732 8094 32734 8146
rect 32786 8094 32788 8146
rect 32732 8036 32788 8094
rect 32732 7970 32788 7980
rect 33068 8148 33124 8158
rect 33068 7812 33124 8092
rect 33180 8036 33236 8046
rect 33180 7942 33236 7980
rect 33404 8036 33460 8046
rect 33404 8034 33572 8036
rect 33404 7982 33406 8034
rect 33458 7982 33572 8034
rect 33404 7980 33572 7982
rect 33404 7970 33460 7980
rect 33068 7756 33460 7812
rect 33404 7586 33460 7756
rect 33404 7534 33406 7586
rect 33458 7534 33460 7586
rect 33404 7522 33460 7534
rect 33516 7588 33572 7980
rect 33516 7522 33572 7532
rect 32060 6690 32228 6692
rect 32060 6638 32062 6690
rect 32114 6638 32228 6690
rect 32060 6636 32228 6638
rect 32508 6972 32676 7028
rect 32060 6626 32116 6636
rect 32508 6580 32564 6972
rect 32620 6804 32676 6814
rect 32620 6690 32676 6748
rect 32956 6692 33012 6702
rect 32620 6638 32622 6690
rect 32674 6638 32676 6690
rect 32620 6626 32676 6638
rect 32844 6636 32956 6692
rect 32508 6514 32564 6524
rect 31500 6466 31556 6478
rect 31500 6414 31502 6466
rect 31554 6414 31556 6466
rect 31500 6018 31556 6414
rect 32172 6356 32228 6366
rect 31500 5966 31502 6018
rect 31554 5966 31556 6018
rect 31500 5954 31556 5966
rect 31612 6018 31668 6030
rect 31612 5966 31614 6018
rect 31666 5966 31668 6018
rect 31612 5236 31668 5966
rect 31612 5170 31668 5180
rect 31836 5906 31892 5918
rect 31836 5854 31838 5906
rect 31890 5854 31892 5906
rect 31836 5010 31892 5854
rect 32172 5122 32228 6300
rect 32732 5236 32788 5246
rect 32732 5142 32788 5180
rect 32172 5070 32174 5122
rect 32226 5070 32228 5122
rect 32172 5058 32228 5070
rect 32844 5122 32900 6636
rect 32956 6626 33012 6636
rect 32844 5070 32846 5122
rect 32898 5070 32900 5122
rect 32844 5058 32900 5070
rect 33180 5012 33236 5022
rect 31836 4958 31838 5010
rect 31890 4958 31892 5010
rect 31836 4946 31892 4958
rect 32956 5010 33460 5012
rect 32956 4958 33182 5010
rect 33234 4958 33460 5010
rect 32956 4956 33460 4958
rect 30828 4510 30830 4562
rect 30882 4510 30884 4562
rect 30604 4340 30660 4350
rect 30604 4246 30660 4284
rect 30828 4228 30884 4510
rect 32284 4900 32340 4910
rect 32284 4450 32340 4844
rect 32284 4398 32286 4450
rect 32338 4398 32340 4450
rect 32284 4386 32340 4398
rect 31836 4340 31892 4350
rect 31388 4228 31444 4238
rect 30828 4226 31444 4228
rect 30828 4174 31390 4226
rect 31442 4174 31444 4226
rect 30828 4172 31444 4174
rect 31388 4162 31444 4172
rect 31836 3556 31892 4284
rect 32956 3666 33012 4956
rect 33180 4946 33236 4956
rect 33068 4564 33124 4574
rect 33068 4470 33124 4508
rect 33404 4338 33460 4956
rect 33628 4452 33684 9324
rect 33964 7474 34020 15148
rect 34076 11396 34132 15484
rect 34412 15314 34468 16156
rect 34412 15262 34414 15314
rect 34466 15262 34468 15314
rect 34412 15250 34468 15262
rect 34524 15316 34580 17052
rect 34636 15986 34692 15998
rect 34636 15934 34638 15986
rect 34690 15934 34692 15986
rect 34636 15540 34692 15934
rect 34860 15986 34916 18060
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35420 17780 35476 17790
rect 35420 16882 35476 17724
rect 35532 17668 35588 18396
rect 35756 18338 35812 18350
rect 35756 18286 35758 18338
rect 35810 18286 35812 18338
rect 35756 17892 35812 18286
rect 35756 17826 35812 17836
rect 35980 17780 36036 19740
rect 36540 20020 36596 20030
rect 36428 19234 36484 19246
rect 36428 19182 36430 19234
rect 36482 19182 36484 19234
rect 36428 18900 36484 19182
rect 36428 18834 36484 18844
rect 36540 18452 36596 19964
rect 36204 18450 36596 18452
rect 36204 18398 36542 18450
rect 36594 18398 36596 18450
rect 36204 18396 36596 18398
rect 35980 17714 36036 17724
rect 36092 18226 36148 18238
rect 36092 18174 36094 18226
rect 36146 18174 36148 18226
rect 35532 17602 35588 17612
rect 35756 17556 35812 17566
rect 35756 17554 36036 17556
rect 35756 17502 35758 17554
rect 35810 17502 36036 17554
rect 35756 17500 36036 17502
rect 35756 17490 35812 17500
rect 35420 16830 35422 16882
rect 35474 16830 35476 16882
rect 35420 16818 35476 16830
rect 35532 16770 35588 16782
rect 35532 16718 35534 16770
rect 35586 16718 35588 16770
rect 34860 15934 34862 15986
rect 34914 15934 34916 15986
rect 34860 15922 34916 15934
rect 35084 16658 35140 16670
rect 35084 16606 35086 16658
rect 35138 16606 35140 16658
rect 35084 15540 35140 16606
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35532 16324 35588 16718
rect 35980 16436 36036 17500
rect 36092 16996 36148 18174
rect 36204 17666 36260 18396
rect 36540 18386 36596 18396
rect 36204 17614 36206 17666
rect 36258 17614 36260 17666
rect 36204 17602 36260 17614
rect 36092 16882 36148 16940
rect 36092 16830 36094 16882
rect 36146 16830 36148 16882
rect 36092 16818 36148 16830
rect 36428 16884 36484 16894
rect 36428 16790 36484 16828
rect 36316 16660 36372 16670
rect 35980 16380 36148 16436
rect 35532 16268 36036 16324
rect 35980 16212 36036 16268
rect 35980 16118 36036 16156
rect 35196 16100 35252 16110
rect 35196 15874 35252 16044
rect 35756 15988 35812 15998
rect 35756 15894 35812 15932
rect 35196 15822 35198 15874
rect 35250 15822 35252 15874
rect 35196 15810 35252 15822
rect 34636 15484 35028 15540
rect 34748 15316 34804 15326
rect 34524 15314 34804 15316
rect 34524 15262 34750 15314
rect 34802 15262 34804 15314
rect 34524 15260 34804 15262
rect 34524 15148 34580 15260
rect 34748 15250 34804 15260
rect 34972 15202 35028 15484
rect 35084 15474 35140 15484
rect 35308 15426 35364 15438
rect 35308 15374 35310 15426
rect 35362 15374 35364 15426
rect 34972 15150 34974 15202
rect 35026 15150 35028 15202
rect 34524 15092 34692 15148
rect 34972 15138 35028 15150
rect 35084 15314 35140 15326
rect 35084 15262 35086 15314
rect 35138 15262 35140 15314
rect 34636 14530 34692 15092
rect 35084 14756 35140 15262
rect 35308 15148 35364 15374
rect 36092 15316 36148 16380
rect 36092 15250 36148 15260
rect 36316 15148 36372 16604
rect 35308 15092 35588 15148
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35532 14756 35588 15092
rect 34636 14478 34638 14530
rect 34690 14478 34692 14530
rect 34636 13636 34692 14478
rect 34972 14700 35140 14756
rect 35196 14700 35588 14756
rect 34972 14420 35028 14700
rect 35084 14532 35140 14542
rect 35084 14438 35140 14476
rect 34972 13746 35028 14364
rect 35084 13860 35140 13870
rect 35084 13766 35140 13804
rect 34972 13694 34974 13746
rect 35026 13694 35028 13746
rect 34972 13682 35028 13694
rect 35196 13748 35252 14700
rect 35532 14644 35588 14700
rect 35532 14578 35588 14588
rect 36204 15092 36372 15148
rect 35308 14530 35364 14542
rect 35308 14478 35310 14530
rect 35362 14478 35364 14530
rect 35308 14308 35364 14478
rect 35756 14308 35812 14318
rect 35308 14306 35812 14308
rect 35308 14254 35758 14306
rect 35810 14254 35812 14306
rect 35308 14252 35812 14254
rect 35308 14196 35364 14252
rect 35756 14242 35812 14252
rect 35308 14130 35364 14140
rect 35196 13682 35252 13692
rect 34636 13542 34692 13580
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 36204 12852 36260 15092
rect 36316 14644 36372 14654
rect 36316 14550 36372 14588
rect 36316 12852 36372 12862
rect 36204 12850 36372 12852
rect 36204 12798 36318 12850
rect 36370 12798 36372 12850
rect 36204 12796 36372 12798
rect 36316 12786 36372 12796
rect 36428 12850 36484 12862
rect 36428 12798 36430 12850
rect 36482 12798 36484 12850
rect 35868 12740 35924 12750
rect 36092 12740 36148 12750
rect 35756 12738 35924 12740
rect 35756 12686 35870 12738
rect 35922 12686 35924 12738
rect 35756 12684 35924 12686
rect 35196 12404 35252 12414
rect 35196 12310 35252 12348
rect 35756 12404 35812 12684
rect 35868 12674 35924 12684
rect 35980 12738 36148 12740
rect 35980 12686 36094 12738
rect 36146 12686 36148 12738
rect 35980 12684 36148 12686
rect 35980 12404 36036 12684
rect 36092 12674 36148 12684
rect 35756 12338 35812 12348
rect 35868 12348 36036 12404
rect 36428 12404 36484 12798
rect 35868 12290 35924 12348
rect 36428 12338 36484 12348
rect 35868 12238 35870 12290
rect 35922 12238 35924 12290
rect 35868 12226 35924 12238
rect 34748 12180 34804 12190
rect 34748 12086 34804 12124
rect 35980 12180 36036 12190
rect 35980 12086 36036 12124
rect 35868 11956 35924 11966
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 34076 11302 34132 11340
rect 34188 11620 34244 11630
rect 34188 10722 34244 11564
rect 34188 10670 34190 10722
rect 34242 10670 34244 10722
rect 34076 10388 34132 10398
rect 34076 9826 34132 10332
rect 34076 9774 34078 9826
rect 34130 9774 34132 9826
rect 34076 9762 34132 9774
rect 34188 9716 34244 10670
rect 34300 11508 34356 11518
rect 34300 10050 34356 11452
rect 34748 11508 34804 11518
rect 34636 11396 34692 11406
rect 34524 11284 34580 11294
rect 34524 11190 34580 11228
rect 34300 9998 34302 10050
rect 34354 9998 34356 10050
rect 34300 9986 34356 9998
rect 34636 10050 34692 11340
rect 34748 11394 34804 11452
rect 34748 11342 34750 11394
rect 34802 11342 34804 11394
rect 34748 11330 34804 11342
rect 35196 11508 35252 11518
rect 35196 11394 35252 11452
rect 35196 11342 35198 11394
rect 35250 11342 35252 11394
rect 35196 11330 35252 11342
rect 35308 11396 35364 11406
rect 35308 11302 35364 11340
rect 34972 11170 35028 11182
rect 34972 11118 34974 11170
rect 35026 11118 35028 11170
rect 34972 10948 35028 11118
rect 34748 10892 35028 10948
rect 34748 10834 34804 10892
rect 34748 10782 34750 10834
rect 34802 10782 34804 10834
rect 34748 10770 34804 10782
rect 34972 10724 35028 10734
rect 34972 10630 35028 10668
rect 35420 10610 35476 10622
rect 35420 10558 35422 10610
rect 35474 10558 35476 10610
rect 34860 10500 34916 10510
rect 34636 9998 34638 10050
rect 34690 9998 34692 10050
rect 34636 9986 34692 9998
rect 34748 10498 34916 10500
rect 34748 10446 34862 10498
rect 34914 10446 34916 10498
rect 34748 10444 34916 10446
rect 34524 9716 34580 9726
rect 34188 9714 34580 9716
rect 34188 9662 34526 9714
rect 34578 9662 34580 9714
rect 34188 9660 34580 9662
rect 34524 9650 34580 9660
rect 34412 7588 34468 7598
rect 34412 7494 34468 7532
rect 33964 7422 33966 7474
rect 34018 7422 34020 7474
rect 33964 6692 34020 7422
rect 33964 6598 34020 6636
rect 34636 7362 34692 7374
rect 34636 7310 34638 7362
rect 34690 7310 34692 7362
rect 34636 5348 34692 7310
rect 34748 6916 34804 10444
rect 34860 10434 34916 10444
rect 35420 10388 35476 10558
rect 35868 10388 35924 11900
rect 36092 11732 36148 11742
rect 36092 11508 36148 11676
rect 36652 11620 36708 20132
rect 37100 19906 37156 26796
rect 37212 26786 37268 26796
rect 37324 26516 37380 28590
rect 37548 28644 37604 28654
rect 37436 27636 37492 27646
rect 37436 26962 37492 27580
rect 37436 26910 37438 26962
rect 37490 26910 37492 26962
rect 37436 26898 37492 26910
rect 37212 26460 37380 26516
rect 37212 24612 37268 26460
rect 37548 26404 37604 28588
rect 37772 28642 37828 28654
rect 37772 28590 37774 28642
rect 37826 28590 37828 28642
rect 37772 27636 37828 28590
rect 38220 28644 38276 28654
rect 38220 28550 38276 28588
rect 38332 28532 38388 29486
rect 38332 28308 38388 28476
rect 38556 28530 38612 29932
rect 39228 29988 39284 29998
rect 39228 29894 39284 29932
rect 39564 29986 39620 29998
rect 39564 29934 39566 29986
rect 39618 29934 39620 29986
rect 39452 29652 39508 29662
rect 38556 28478 38558 28530
rect 38610 28478 38612 28530
rect 38556 28466 38612 28478
rect 38780 29538 38836 29550
rect 38780 29486 38782 29538
rect 38834 29486 38836 29538
rect 38780 28420 38836 29486
rect 39116 29426 39172 29438
rect 39116 29374 39118 29426
rect 39170 29374 39172 29426
rect 39116 29316 39172 29374
rect 39452 29426 39508 29596
rect 39452 29374 39454 29426
rect 39506 29374 39508 29426
rect 39452 29362 39508 29374
rect 39116 29250 39172 29260
rect 39564 29316 39620 29934
rect 42700 29426 42756 30942
rect 43036 31892 43092 31902
rect 43036 30994 43092 31836
rect 43036 30942 43038 30994
rect 43090 30942 43092 30994
rect 43036 30930 43092 30942
rect 42700 29374 42702 29426
rect 42754 29374 42756 29426
rect 42700 29362 42756 29374
rect 43260 29428 43316 29438
rect 43260 29334 43316 29372
rect 39564 29250 39620 29260
rect 40236 29316 40292 29326
rect 38780 28354 38836 28364
rect 39788 29202 39844 29214
rect 39788 29150 39790 29202
rect 39842 29150 39844 29202
rect 39788 28420 39844 29150
rect 38332 28252 38724 28308
rect 38220 27972 38276 27982
rect 38556 27972 38612 27982
rect 38220 27970 38612 27972
rect 38220 27918 38222 27970
rect 38274 27918 38558 27970
rect 38610 27918 38612 27970
rect 38220 27916 38612 27918
rect 38220 27906 38276 27916
rect 38556 27906 38612 27916
rect 38668 27970 38724 28252
rect 38668 27918 38670 27970
rect 38722 27918 38724 27970
rect 38668 27906 38724 27918
rect 39788 27860 39844 28364
rect 39788 27794 39844 27804
rect 38556 27636 38612 27646
rect 37772 27634 38612 27636
rect 37772 27582 38558 27634
rect 38610 27582 38612 27634
rect 37772 27580 38612 27582
rect 37324 26348 37604 26404
rect 37324 25394 37380 26348
rect 37324 25342 37326 25394
rect 37378 25342 37380 25394
rect 37324 24948 37380 25342
rect 37996 25506 38052 25518
rect 37996 25454 37998 25506
rect 38050 25454 38052 25506
rect 37324 24882 37380 24892
rect 37884 25284 37940 25294
rect 37884 24722 37940 25228
rect 37884 24670 37886 24722
rect 37938 24670 37940 24722
rect 37884 24658 37940 24670
rect 37324 24612 37380 24622
rect 37996 24612 38052 25454
rect 38556 25506 38612 27580
rect 38780 27074 38836 27086
rect 38780 27022 38782 27074
rect 38834 27022 38836 27074
rect 38780 26908 38836 27022
rect 39228 27076 39284 27086
rect 39228 26982 39284 27020
rect 40236 26908 40292 29260
rect 42588 28084 42644 28094
rect 41356 27972 41412 27982
rect 40796 27860 40852 27870
rect 40796 27766 40852 27804
rect 41356 27858 41412 27916
rect 41356 27806 41358 27858
rect 41410 27806 41412 27858
rect 38780 26852 39060 26908
rect 39004 26404 39060 26852
rect 39676 26852 40292 26908
rect 39676 26516 39732 26852
rect 39788 26516 39844 26526
rect 39340 26514 39844 26516
rect 39340 26462 39790 26514
rect 39842 26462 39844 26514
rect 39340 26460 39844 26462
rect 39228 26404 39284 26414
rect 39004 26402 39284 26404
rect 39004 26350 39230 26402
rect 39282 26350 39284 26402
rect 39004 26348 39284 26350
rect 38892 26290 38948 26302
rect 38892 26238 38894 26290
rect 38946 26238 38948 26290
rect 38892 26068 38948 26238
rect 39228 26292 39284 26348
rect 39228 26226 39284 26236
rect 39340 26068 39396 26460
rect 39788 26450 39844 26460
rect 38892 26012 39396 26068
rect 38556 25454 38558 25506
rect 38610 25454 38612 25506
rect 38556 25442 38612 25454
rect 38668 25394 38724 25406
rect 38668 25342 38670 25394
rect 38722 25342 38724 25394
rect 38668 24836 38724 25342
rect 38892 24948 38948 24958
rect 38892 24854 38948 24892
rect 38780 24836 38836 24846
rect 38108 24834 38836 24836
rect 38108 24782 38782 24834
rect 38834 24782 38836 24834
rect 38108 24780 38836 24782
rect 38108 24722 38164 24780
rect 38780 24770 38836 24780
rect 41356 24836 41412 27806
rect 41468 27188 41524 27198
rect 41468 26962 41524 27132
rect 42588 27188 42644 28028
rect 42588 27094 42644 27132
rect 41468 26910 41470 26962
rect 41522 26910 41524 26962
rect 41468 26898 41524 26910
rect 42364 27076 42420 27086
rect 42252 26852 42308 26862
rect 41356 24742 41412 24780
rect 41804 26850 42308 26852
rect 41804 26798 42254 26850
rect 42306 26798 42308 26850
rect 41804 26796 42308 26798
rect 38108 24670 38110 24722
rect 38162 24670 38164 24722
rect 38108 24658 38164 24670
rect 39116 24724 39172 24734
rect 39116 24722 40068 24724
rect 39116 24670 39118 24722
rect 39170 24670 40068 24722
rect 39116 24668 40068 24670
rect 39116 24658 39172 24668
rect 37212 24610 37604 24612
rect 37212 24558 37326 24610
rect 37378 24558 37604 24610
rect 37212 24556 37604 24558
rect 37324 24546 37380 24556
rect 37212 23380 37268 23390
rect 37212 22258 37268 23324
rect 37212 22206 37214 22258
rect 37266 22206 37268 22258
rect 37212 22194 37268 22206
rect 37324 22258 37380 22270
rect 37324 22206 37326 22258
rect 37378 22206 37380 22258
rect 37324 21924 37380 22206
rect 37436 22260 37492 22270
rect 37548 22260 37604 24556
rect 37996 24546 38052 24556
rect 38444 24500 38500 24510
rect 38444 24498 38612 24500
rect 38444 24446 38446 24498
rect 38498 24446 38612 24498
rect 38444 24444 38612 24446
rect 38444 24434 38500 24444
rect 38444 23380 38500 23390
rect 38332 23044 38388 23054
rect 37772 22484 37828 22494
rect 37772 22390 37828 22428
rect 38332 22482 38388 22988
rect 38332 22430 38334 22482
rect 38386 22430 38388 22482
rect 38332 22418 38388 22430
rect 38444 22260 38500 23324
rect 38556 22372 38612 24444
rect 38892 23156 38948 23166
rect 38948 23100 39060 23156
rect 38892 23062 38948 23100
rect 38556 22316 38948 22372
rect 37548 22204 37828 22260
rect 38444 22204 38836 22260
rect 37436 22166 37492 22204
rect 37324 21858 37380 21868
rect 37548 21700 37604 21710
rect 37548 21698 37716 21700
rect 37548 21646 37550 21698
rect 37602 21646 37716 21698
rect 37548 21644 37716 21646
rect 37548 21634 37604 21644
rect 37660 20914 37716 21644
rect 37660 20862 37662 20914
rect 37714 20862 37716 20914
rect 37100 19854 37102 19906
rect 37154 19854 37156 19906
rect 37100 19124 37156 19854
rect 37436 19908 37492 19918
rect 37436 19234 37492 19852
rect 37660 19796 37716 20862
rect 37660 19730 37716 19740
rect 37436 19182 37438 19234
rect 37490 19182 37492 19234
rect 37212 19124 37268 19134
rect 37100 19122 37268 19124
rect 37100 19070 37214 19122
rect 37266 19070 37268 19122
rect 37100 19068 37268 19070
rect 37100 18452 37156 19068
rect 37212 19058 37268 19068
rect 36988 18226 37044 18238
rect 36988 18174 36990 18226
rect 37042 18174 37044 18226
rect 36988 17892 37044 18174
rect 36988 17826 37044 17836
rect 36988 17220 37044 17230
rect 36764 16884 36820 16894
rect 36764 16790 36820 16828
rect 36988 15148 37044 17164
rect 37100 15986 37156 18396
rect 37212 18900 37268 18910
rect 37212 18450 37268 18844
rect 37436 18564 37492 19182
rect 37772 18676 37828 22204
rect 38556 22036 38612 22046
rect 38556 21588 38612 21980
rect 38668 21588 38724 21598
rect 38612 21586 38724 21588
rect 38612 21534 38670 21586
rect 38722 21534 38724 21586
rect 38612 21532 38724 21534
rect 38556 21494 38612 21532
rect 38668 21522 38724 21532
rect 38108 21028 38164 21038
rect 38108 20802 38164 20972
rect 38668 21028 38724 21038
rect 38668 20914 38724 20972
rect 38668 20862 38670 20914
rect 38722 20862 38724 20914
rect 38668 20850 38724 20862
rect 38108 20750 38110 20802
rect 38162 20750 38164 20802
rect 38108 20738 38164 20750
rect 38780 20188 38836 22204
rect 37884 20132 37940 20142
rect 37884 20018 37940 20076
rect 38668 20132 38836 20188
rect 37884 19966 37886 20018
rect 37938 19966 37940 20018
rect 37884 19954 37940 19966
rect 38332 20018 38388 20030
rect 38332 19966 38334 20018
rect 38386 19966 38388 20018
rect 38332 19796 38388 19966
rect 38556 20018 38612 20030
rect 38556 19966 38558 20018
rect 38610 19966 38612 20018
rect 38332 19730 38388 19740
rect 38444 19906 38500 19918
rect 38444 19854 38446 19906
rect 38498 19854 38500 19906
rect 37660 18620 37828 18676
rect 38220 19346 38276 19358
rect 38220 19294 38222 19346
rect 38274 19294 38276 19346
rect 37548 18564 37604 18574
rect 37436 18562 37604 18564
rect 37436 18510 37550 18562
rect 37602 18510 37604 18562
rect 37436 18508 37604 18510
rect 37548 18498 37604 18508
rect 37212 18398 37214 18450
rect 37266 18398 37268 18450
rect 37212 18386 37268 18398
rect 37436 18340 37492 18350
rect 37324 18338 37492 18340
rect 37324 18286 37438 18338
rect 37490 18286 37492 18338
rect 37324 18284 37492 18286
rect 37100 15934 37102 15986
rect 37154 15934 37156 15986
rect 37100 15922 37156 15934
rect 37212 17444 37268 17454
rect 37212 16884 37268 17388
rect 37212 15314 37268 16828
rect 37212 15262 37214 15314
rect 37266 15262 37268 15314
rect 37212 15250 37268 15262
rect 36988 15092 37156 15148
rect 36988 13634 37044 13646
rect 36988 13582 36990 13634
rect 37042 13582 37044 13634
rect 36876 12404 36932 12414
rect 36876 12178 36932 12348
rect 36876 12126 36878 12178
rect 36930 12126 36932 12178
rect 36876 12114 36932 12126
rect 36876 11954 36932 11966
rect 36876 11902 36878 11954
rect 36930 11902 36932 11954
rect 36876 11620 36932 11902
rect 36988 11844 37044 13582
rect 36988 11778 37044 11788
rect 36876 11564 37044 11620
rect 36652 11554 36708 11564
rect 36092 10834 36148 11452
rect 36876 11396 36932 11406
rect 36092 10782 36094 10834
rect 36146 10782 36148 10834
rect 36092 10770 36148 10782
rect 36316 11394 36932 11396
rect 36316 11342 36878 11394
rect 36930 11342 36932 11394
rect 36316 11340 36932 11342
rect 36316 10834 36372 11340
rect 36876 11330 36932 11340
rect 36988 11172 37044 11564
rect 36316 10782 36318 10834
rect 36370 10782 36372 10834
rect 36316 10770 36372 10782
rect 36876 11116 37044 11172
rect 35980 10612 36036 10622
rect 35980 10518 36036 10556
rect 35868 10332 36036 10388
rect 35420 10322 35476 10332
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35868 9940 35924 9950
rect 35868 9846 35924 9884
rect 35756 9604 35812 9614
rect 35308 9602 35812 9604
rect 35308 9550 35758 9602
rect 35810 9550 35812 9602
rect 35308 9548 35812 9550
rect 35308 9042 35364 9548
rect 35308 8990 35310 9042
rect 35362 8990 35364 9042
rect 35308 8978 35364 8990
rect 34972 8818 35028 8830
rect 34972 8766 34974 8818
rect 35026 8766 35028 8818
rect 34860 7700 34916 7710
rect 34860 7474 34916 7644
rect 34860 7422 34862 7474
rect 34914 7422 34916 7474
rect 34860 7410 34916 7422
rect 34748 6860 34916 6916
rect 34748 5348 34804 5358
rect 33964 5346 34804 5348
rect 33964 5294 34750 5346
rect 34802 5294 34804 5346
rect 33964 5292 34804 5294
rect 33964 5122 34020 5292
rect 34748 5282 34804 5292
rect 33964 5070 33966 5122
rect 34018 5070 34020 5122
rect 33964 5058 34020 5070
rect 34076 5180 34580 5236
rect 34076 5010 34132 5180
rect 34524 5124 34580 5180
rect 34860 5124 34916 6860
rect 34524 5122 34916 5124
rect 34524 5070 34526 5122
rect 34578 5070 34916 5122
rect 34524 5068 34916 5070
rect 34524 5058 34580 5068
rect 34076 4958 34078 5010
rect 34130 4958 34132 5010
rect 34076 4946 34132 4958
rect 34300 5012 34356 5022
rect 34300 4918 34356 4956
rect 34076 4564 34132 4574
rect 34076 4470 34132 4508
rect 33404 4286 33406 4338
rect 33458 4286 33460 4338
rect 33404 4274 33460 4286
rect 33516 4450 33684 4452
rect 33516 4398 33630 4450
rect 33682 4398 33684 4450
rect 33516 4396 33684 4398
rect 33516 4116 33572 4396
rect 33628 4386 33684 4396
rect 34524 4452 34580 4462
rect 34524 4358 34580 4396
rect 34300 4340 34356 4350
rect 34300 4246 34356 4284
rect 34972 4340 35028 8766
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35308 8372 35364 8382
rect 35308 8278 35364 8316
rect 35532 8258 35588 9548
rect 35756 9538 35812 9548
rect 35980 9042 36036 10332
rect 36092 9268 36148 9278
rect 36092 9154 36148 9212
rect 36764 9268 36820 9278
rect 36764 9174 36820 9212
rect 36092 9102 36094 9154
rect 36146 9102 36148 9154
rect 36092 9090 36148 9102
rect 35980 8990 35982 9042
rect 36034 8990 36036 9042
rect 35980 8978 36036 8990
rect 35532 8206 35534 8258
rect 35586 8206 35588 8258
rect 35532 8194 35588 8206
rect 36092 8148 36148 8158
rect 36092 8054 36148 8092
rect 35532 8036 35588 8046
rect 35532 7698 35588 7980
rect 35532 7646 35534 7698
rect 35586 7646 35588 7698
rect 35532 7634 35588 7646
rect 36092 7700 36148 7710
rect 36092 7606 36148 7644
rect 35308 7474 35364 7486
rect 35308 7422 35310 7474
rect 35362 7422 35364 7474
rect 35308 7364 35364 7422
rect 35084 7308 35364 7364
rect 35644 7474 35700 7486
rect 35644 7422 35646 7474
rect 35698 7422 35700 7474
rect 35084 6578 35140 7308
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35644 6804 35700 7422
rect 35644 6738 35700 6748
rect 35868 6914 35924 6926
rect 35868 6862 35870 6914
rect 35922 6862 35924 6914
rect 35084 6526 35086 6578
rect 35138 6526 35140 6578
rect 35084 6514 35140 6526
rect 35196 6690 35252 6702
rect 35196 6638 35198 6690
rect 35250 6638 35252 6690
rect 35196 6356 35252 6638
rect 35196 6290 35252 6300
rect 35868 6692 35924 6862
rect 35868 6018 35924 6636
rect 35868 5966 35870 6018
rect 35922 5966 35924 6018
rect 35868 5954 35924 5966
rect 36876 6692 36932 11116
rect 37100 9268 37156 15092
rect 37324 13746 37380 18284
rect 37436 18274 37492 18284
rect 37660 17220 37716 18620
rect 37772 18452 37828 18462
rect 37772 18358 37828 18396
rect 38220 17444 38276 19294
rect 38332 19236 38388 19246
rect 38332 19142 38388 19180
rect 38444 18452 38500 19854
rect 38556 19348 38612 19966
rect 38556 19282 38612 19292
rect 38556 19122 38612 19134
rect 38556 19070 38558 19122
rect 38610 19070 38612 19122
rect 38556 18564 38612 19070
rect 38556 18498 38612 18508
rect 38444 18386 38500 18396
rect 38556 18340 38612 18350
rect 38556 18246 38612 18284
rect 38444 18226 38500 18238
rect 38444 18174 38446 18226
rect 38498 18174 38500 18226
rect 38444 17892 38500 18174
rect 38444 17826 38500 17836
rect 38332 17444 38388 17454
rect 38220 17388 38332 17444
rect 38332 17378 38388 17388
rect 37660 17154 37716 17164
rect 37660 16996 37716 17006
rect 37716 16940 37828 16996
rect 37660 16902 37716 16940
rect 37548 16884 37604 16894
rect 37436 16882 37604 16884
rect 37436 16830 37550 16882
rect 37602 16830 37604 16882
rect 37436 16828 37604 16830
rect 37436 16212 37492 16828
rect 37548 16818 37604 16828
rect 37772 16324 37828 16940
rect 37884 16772 37940 16782
rect 37884 16770 38052 16772
rect 37884 16718 37886 16770
rect 37938 16718 38052 16770
rect 37884 16716 38052 16718
rect 37884 16706 37940 16716
rect 37884 16324 37940 16334
rect 37772 16322 37940 16324
rect 37772 16270 37886 16322
rect 37938 16270 37940 16322
rect 37772 16268 37940 16270
rect 37884 16258 37940 16268
rect 37436 16098 37492 16156
rect 37436 16046 37438 16098
rect 37490 16046 37492 16098
rect 37436 16034 37492 16046
rect 37996 16100 38052 16716
rect 37996 16044 38388 16100
rect 38220 15876 38276 15886
rect 38220 15782 38276 15820
rect 37436 15316 37492 15326
rect 37436 15222 37492 15260
rect 37772 15316 37828 15326
rect 38108 15316 38164 15326
rect 37772 15314 38164 15316
rect 37772 15262 37774 15314
rect 37826 15262 38110 15314
rect 38162 15262 38164 15314
rect 37772 15260 38164 15262
rect 37772 15250 37828 15260
rect 37884 14530 37940 15260
rect 38108 15250 38164 15260
rect 38220 15316 38276 15326
rect 38220 15148 38276 15260
rect 38332 15314 38388 16044
rect 38668 16098 38724 20132
rect 38668 16046 38670 16098
rect 38722 16046 38724 16098
rect 38668 16034 38724 16046
rect 38780 18452 38836 18462
rect 38892 18452 38948 22316
rect 39004 22370 39060 23100
rect 39116 23044 39172 23054
rect 39172 22988 39284 23044
rect 39116 22950 39172 22988
rect 39228 22482 39284 22988
rect 39228 22430 39230 22482
rect 39282 22430 39284 22482
rect 39228 22418 39284 22430
rect 39340 22930 39396 22942
rect 39340 22878 39342 22930
rect 39394 22878 39396 22930
rect 39004 22318 39006 22370
rect 39058 22318 39060 22370
rect 39004 22306 39060 22318
rect 39228 21474 39284 21486
rect 39228 21422 39230 21474
rect 39282 21422 39284 21474
rect 39228 20804 39284 21422
rect 39340 21252 39396 22878
rect 40012 22484 40068 24668
rect 40572 24612 40628 24622
rect 39564 22428 40068 22484
rect 39564 21586 39620 22428
rect 40012 22370 40068 22428
rect 40012 22318 40014 22370
rect 40066 22318 40068 22370
rect 40012 22306 40068 22318
rect 40460 22482 40516 22494
rect 40460 22430 40462 22482
rect 40514 22430 40516 22482
rect 39676 22260 39732 22270
rect 39676 22258 39956 22260
rect 39676 22206 39678 22258
rect 39730 22206 39956 22258
rect 39676 22204 39956 22206
rect 39676 22194 39732 22204
rect 39564 21534 39566 21586
rect 39618 21534 39620 21586
rect 39564 21522 39620 21534
rect 39900 21252 39956 22204
rect 39900 21196 40068 21252
rect 39340 21186 39396 21196
rect 39676 20804 39732 20814
rect 39228 20802 39732 20804
rect 39228 20750 39678 20802
rect 39730 20750 39732 20802
rect 39228 20748 39732 20750
rect 39228 20188 39284 20748
rect 39676 20738 39732 20748
rect 38780 18450 38948 18452
rect 38780 18398 38782 18450
rect 38834 18398 38948 18450
rect 38780 18396 38948 18398
rect 39004 20132 39284 20188
rect 39900 20690 39956 20702
rect 39900 20638 39902 20690
rect 39954 20638 39956 20690
rect 39452 20132 39508 20142
rect 39900 20132 39956 20638
rect 38780 17442 38836 18396
rect 38780 17390 38782 17442
rect 38834 17390 38836 17442
rect 38332 15262 38334 15314
rect 38386 15262 38388 15314
rect 38332 15250 38388 15262
rect 38220 15092 38388 15148
rect 37884 14478 37886 14530
rect 37938 14478 37940 14530
rect 37884 14466 37940 14478
rect 37772 13860 37828 13870
rect 37772 13766 37828 13804
rect 37324 13694 37326 13746
rect 37378 13694 37380 13746
rect 37324 13682 37380 13694
rect 37996 13748 38052 13758
rect 37212 12066 37268 12078
rect 37212 12014 37214 12066
rect 37266 12014 37268 12066
rect 37212 10612 37268 12014
rect 37324 11620 37380 11630
rect 37324 11394 37380 11564
rect 37436 11508 37492 11518
rect 37436 11506 37940 11508
rect 37436 11454 37438 11506
rect 37490 11454 37940 11506
rect 37436 11452 37940 11454
rect 37436 11442 37492 11452
rect 37324 11342 37326 11394
rect 37378 11342 37380 11394
rect 37324 11330 37380 11342
rect 37884 11394 37940 11452
rect 37884 11342 37886 11394
rect 37938 11342 37940 11394
rect 37884 11330 37940 11342
rect 37996 11282 38052 13692
rect 38332 12404 38388 15092
rect 38556 14980 38612 14990
rect 38444 14924 38556 14980
rect 38444 13858 38500 14924
rect 38556 14914 38612 14924
rect 38556 14644 38612 14654
rect 38556 14550 38612 14588
rect 38444 13806 38446 13858
rect 38498 13806 38500 13858
rect 38444 13524 38500 13806
rect 38668 14420 38724 14430
rect 38668 13858 38724 14364
rect 38668 13806 38670 13858
rect 38722 13806 38724 13858
rect 38668 13748 38724 13806
rect 38668 13682 38724 13692
rect 38780 13636 38836 17390
rect 39004 16100 39060 20132
rect 39452 20130 39956 20132
rect 39452 20078 39454 20130
rect 39506 20078 39956 20130
rect 39452 20076 39956 20078
rect 39340 20020 39396 20030
rect 39340 19926 39396 19964
rect 39452 18900 39508 20076
rect 40012 19908 40068 21196
rect 40236 20804 40292 20814
rect 40236 20242 40292 20748
rect 40236 20190 40238 20242
rect 40290 20190 40292 20242
rect 40236 20178 40292 20190
rect 40348 20690 40404 20702
rect 40348 20638 40350 20690
rect 40402 20638 40404 20690
rect 40012 19842 40068 19852
rect 40124 20132 40180 20142
rect 40124 20020 40180 20076
rect 40348 20020 40404 20638
rect 40124 20018 40404 20020
rect 40124 19966 40126 20018
rect 40178 19966 40404 20018
rect 40124 19964 40404 19966
rect 40460 20020 40516 22430
rect 40124 19684 40180 19964
rect 40012 19628 40180 19684
rect 40012 19234 40068 19628
rect 40012 19182 40014 19234
rect 40066 19182 40068 19234
rect 40012 19170 40068 19182
rect 39452 18834 39508 18844
rect 40124 19122 40180 19134
rect 40124 19070 40126 19122
rect 40178 19070 40180 19122
rect 40124 18900 40180 19070
rect 40236 19124 40292 19134
rect 40460 19124 40516 19964
rect 40236 19122 40516 19124
rect 40236 19070 40238 19122
rect 40290 19070 40516 19122
rect 40236 19068 40516 19070
rect 40236 19058 40292 19068
rect 40124 18834 40180 18844
rect 39228 18452 39284 18462
rect 39228 18358 39284 18396
rect 39452 18450 39508 18462
rect 39452 18398 39454 18450
rect 39506 18398 39508 18450
rect 39340 18340 39396 18350
rect 39452 18340 39508 18398
rect 39396 18284 39508 18340
rect 40124 18340 40180 18350
rect 39340 18274 39396 18284
rect 40124 18246 40180 18284
rect 40348 17556 40404 19068
rect 40572 17668 40628 24556
rect 41692 24612 41748 24622
rect 41692 24518 41748 24556
rect 40796 24108 41300 24164
rect 40796 24050 40852 24108
rect 40796 23998 40798 24050
rect 40850 23998 40852 24050
rect 40796 23986 40852 23998
rect 41132 23938 41188 23950
rect 41132 23886 41134 23938
rect 41186 23886 41188 23938
rect 41132 23828 41188 23886
rect 41244 23940 41300 24108
rect 41692 23940 41748 23950
rect 41804 23940 41860 26796
rect 42252 26786 42308 26796
rect 42252 26292 42308 26302
rect 42252 26198 42308 26236
rect 42364 25620 42420 27020
rect 43036 27076 43092 27086
rect 43372 27076 43428 33068
rect 43484 33058 43540 33068
rect 43596 33236 43652 33246
rect 43596 32674 43652 33180
rect 43708 33012 43764 33294
rect 43708 32946 43764 32956
rect 43596 32622 43598 32674
rect 43650 32622 43652 32674
rect 43596 32610 43652 32622
rect 43708 32788 43764 32798
rect 43820 32788 43876 33516
rect 43708 32786 43876 32788
rect 43708 32734 43710 32786
rect 43762 32734 43876 32786
rect 43708 32732 43876 32734
rect 43708 31892 43764 32732
rect 43932 32676 43988 32686
rect 43932 32582 43988 32620
rect 43708 31826 43764 31836
rect 44044 31780 44100 37436
rect 44268 37378 44324 37390
rect 44268 37326 44270 37378
rect 44322 37326 44324 37378
rect 44156 37266 44212 37278
rect 44156 37214 44158 37266
rect 44210 37214 44212 37266
rect 44156 36708 44212 37214
rect 44268 37044 44324 37326
rect 44268 36978 44324 36988
rect 44156 36642 44212 36652
rect 44380 34356 44436 38612
rect 44492 37268 44548 37278
rect 44492 37174 44548 37212
rect 44492 34356 44548 34366
rect 44380 34354 44548 34356
rect 44380 34302 44494 34354
rect 44546 34302 44548 34354
rect 44380 34300 44548 34302
rect 44492 34290 44548 34300
rect 44604 33572 44660 38612
rect 44716 37266 44772 37278
rect 44716 37214 44718 37266
rect 44770 37214 44772 37266
rect 44716 36708 44772 37214
rect 44828 37044 44884 38612
rect 44940 37268 44996 39900
rect 45164 39620 45220 39630
rect 45276 39620 45332 40350
rect 46284 40404 46340 40908
rect 46284 40310 46340 40348
rect 45164 39618 45332 39620
rect 45164 39566 45166 39618
rect 45218 39566 45332 39618
rect 45164 39564 45332 39566
rect 45836 39618 45892 39630
rect 45836 39566 45838 39618
rect 45890 39566 45892 39618
rect 45164 39554 45220 39564
rect 45612 38948 45668 38958
rect 45836 38948 45892 39566
rect 46060 39620 46116 39630
rect 45668 38892 45892 38948
rect 45948 39506 46004 39518
rect 45948 39454 45950 39506
rect 46002 39454 46004 39506
rect 45948 39060 46004 39454
rect 45612 38854 45668 38892
rect 45052 38834 45108 38846
rect 45052 38782 45054 38834
rect 45106 38782 45108 38834
rect 45052 38164 45108 38782
rect 45164 38836 45220 38846
rect 45164 38742 45220 38780
rect 45948 38834 46004 39004
rect 45948 38782 45950 38834
rect 46002 38782 46004 38834
rect 45948 38770 46004 38782
rect 46060 38274 46116 39564
rect 46284 39396 46340 39406
rect 46284 38946 46340 39340
rect 46284 38894 46286 38946
rect 46338 38894 46340 38946
rect 46284 38882 46340 38894
rect 46396 38836 46452 38846
rect 46396 38742 46452 38780
rect 46508 38668 46564 41916
rect 46620 41860 46676 42140
rect 47516 42084 47572 42094
rect 47516 41990 47572 42028
rect 47292 41972 47348 41982
rect 47292 41878 47348 41916
rect 46620 41804 46900 41860
rect 46732 41636 46788 41646
rect 46620 41300 46676 41310
rect 46620 41206 46676 41244
rect 46732 41074 46788 41580
rect 46732 41022 46734 41074
rect 46786 41022 46788 41074
rect 46732 40964 46788 41022
rect 46732 40898 46788 40908
rect 46732 40404 46788 40414
rect 46844 40404 46900 41804
rect 47068 41746 47124 41758
rect 47068 41694 47070 41746
rect 47122 41694 47124 41746
rect 47068 41412 47124 41694
rect 47068 41346 47124 41356
rect 47292 41748 47348 41758
rect 47292 41410 47348 41692
rect 47292 41358 47294 41410
rect 47346 41358 47348 41410
rect 47292 41346 47348 41358
rect 47516 41188 47572 41198
rect 47628 41188 47684 50372
rect 47740 48802 47796 48814
rect 47740 48750 47742 48802
rect 47794 48750 47796 48802
rect 47740 48132 47796 48750
rect 48412 48356 48468 48366
rect 47740 48038 47796 48076
rect 47964 48244 48020 48254
rect 47852 48020 47908 48030
rect 47852 47926 47908 47964
rect 47852 47684 47908 47694
rect 47964 47684 48020 48188
rect 47852 47682 48020 47684
rect 47852 47630 47854 47682
rect 47906 47630 48020 47682
rect 47852 47628 48020 47630
rect 47852 47618 47908 47628
rect 48076 47346 48132 47358
rect 48076 47294 48078 47346
rect 48130 47294 48132 47346
rect 47964 46004 48020 46014
rect 48076 46004 48132 47294
rect 47964 46002 48076 46004
rect 47964 45950 47966 46002
rect 48018 45950 48076 46002
rect 47964 45948 48076 45950
rect 47964 45938 48020 45948
rect 48076 45910 48132 45948
rect 48412 45666 48468 48300
rect 48412 45614 48414 45666
rect 48466 45614 48468 45666
rect 48412 45332 48468 45614
rect 47740 45220 47796 45230
rect 47740 45126 47796 45164
rect 48412 43764 48468 45276
rect 48412 43698 48468 43708
rect 47740 43540 47796 43550
rect 47740 41970 47796 43484
rect 47964 42754 48020 42766
rect 47964 42702 47966 42754
rect 48018 42702 48020 42754
rect 47740 41918 47742 41970
rect 47794 41918 47796 41970
rect 47740 41906 47796 41918
rect 47852 41972 47908 41982
rect 47852 41878 47908 41916
rect 47516 41186 47628 41188
rect 47516 41134 47518 41186
rect 47570 41134 47628 41186
rect 47516 41132 47628 41134
rect 47516 41122 47572 41132
rect 46732 40402 47012 40404
rect 46732 40350 46734 40402
rect 46786 40350 47012 40402
rect 46732 40348 47012 40350
rect 46732 40338 46788 40348
rect 46732 39618 46788 39630
rect 46732 39566 46734 39618
rect 46786 39566 46788 39618
rect 46060 38222 46062 38274
rect 46114 38222 46116 38274
rect 46060 38210 46116 38222
rect 46172 38612 46564 38668
rect 46620 39396 46676 39406
rect 46732 39396 46788 39566
rect 46676 39340 46788 39396
rect 46844 39396 46900 39406
rect 45276 38164 45332 38174
rect 45052 38162 45332 38164
rect 45052 38110 45278 38162
rect 45330 38110 45332 38162
rect 45052 38108 45332 38110
rect 45052 37492 45108 38108
rect 45276 38098 45332 38108
rect 45052 37426 45108 37436
rect 45388 38050 45444 38062
rect 45388 37998 45390 38050
rect 45442 37998 45444 38050
rect 45276 37268 45332 37278
rect 44940 37266 45332 37268
rect 44940 37214 45278 37266
rect 45330 37214 45332 37266
rect 44940 37212 45332 37214
rect 44940 37044 44996 37054
rect 44828 36988 44940 37044
rect 44940 36820 44996 36988
rect 44940 36764 45108 36820
rect 44716 36642 44772 36652
rect 44828 36482 44884 36494
rect 44828 36430 44830 36482
rect 44882 36430 44884 36482
rect 44828 35476 44884 36430
rect 44828 34914 44884 35420
rect 44940 36372 44996 36382
rect 44940 35138 44996 36316
rect 44940 35086 44942 35138
rect 44994 35086 44996 35138
rect 44940 35074 44996 35086
rect 44828 34862 44830 34914
rect 44882 34862 44884 34914
rect 44828 34850 44884 34862
rect 44940 34804 44996 34814
rect 45052 34804 45108 36764
rect 45276 36484 45332 37212
rect 45388 37044 45444 37998
rect 45724 37268 45780 37278
rect 45948 37268 46004 37278
rect 45724 37174 45780 37212
rect 45836 37212 45948 37268
rect 45388 36978 45444 36988
rect 45276 36418 45332 36428
rect 45724 35698 45780 35710
rect 45724 35646 45726 35698
rect 45778 35646 45780 35698
rect 45724 35588 45780 35646
rect 45724 35522 45780 35532
rect 44940 34802 45108 34804
rect 44940 34750 44942 34802
rect 44994 34750 45108 34802
rect 44940 34748 45108 34750
rect 45164 34804 45220 34814
rect 44940 34738 44996 34748
rect 44604 33506 44660 33516
rect 45164 34130 45220 34748
rect 45388 34244 45444 34254
rect 45388 34242 45556 34244
rect 45388 34190 45390 34242
rect 45442 34190 45556 34242
rect 45388 34188 45556 34190
rect 45388 34178 45444 34188
rect 45164 34078 45166 34130
rect 45218 34078 45220 34130
rect 45164 33458 45220 34078
rect 45164 33406 45166 33458
rect 45218 33406 45220 33458
rect 45164 33394 45220 33406
rect 45388 33684 45444 33694
rect 45276 33348 45332 33358
rect 45276 33254 45332 33292
rect 44044 31714 44100 31724
rect 44156 31892 44212 31902
rect 44156 30098 44212 31836
rect 45388 31220 45444 33628
rect 45500 33236 45556 34188
rect 45612 33236 45668 33246
rect 45500 33180 45612 33236
rect 45612 33170 45668 33180
rect 45388 31126 45444 31164
rect 44156 30046 44158 30098
rect 44210 30046 44212 30098
rect 44156 30034 44212 30046
rect 44268 30100 44324 30110
rect 44268 30006 44324 30044
rect 45612 30100 45668 30110
rect 45612 30006 45668 30044
rect 45836 30098 45892 37212
rect 45948 37174 46004 37212
rect 46060 37154 46116 37166
rect 46060 37102 46062 37154
rect 46114 37102 46116 37154
rect 45948 36706 46004 36718
rect 45948 36654 45950 36706
rect 46002 36654 46004 36706
rect 45948 34130 46004 36654
rect 46060 36708 46116 37102
rect 46060 36642 46116 36652
rect 46060 36484 46116 36494
rect 46060 36390 46116 36428
rect 45948 34078 45950 34130
rect 46002 34078 46004 34130
rect 45948 33348 46004 34078
rect 45948 33282 46004 33292
rect 46172 31890 46228 38612
rect 46620 38500 46676 39340
rect 46844 39302 46900 39340
rect 46284 38444 46676 38500
rect 46284 35698 46340 38444
rect 46956 37268 47012 40348
rect 47292 40292 47348 40302
rect 47292 38834 47348 40236
rect 47292 38782 47294 38834
rect 47346 38782 47348 38834
rect 47292 38770 47348 38782
rect 46956 36596 47012 37212
rect 47180 36708 47236 36718
rect 46956 36540 47124 36596
rect 47068 36482 47124 36540
rect 47068 36430 47070 36482
rect 47122 36430 47124 36482
rect 47068 36418 47124 36430
rect 46284 35646 46286 35698
rect 46338 35646 46340 35698
rect 46284 35634 46340 35646
rect 47180 35698 47236 36652
rect 47292 36372 47348 36382
rect 47292 36278 47348 36316
rect 47180 35646 47182 35698
rect 47234 35646 47236 35698
rect 46732 35588 46788 35598
rect 46732 35476 46788 35532
rect 46732 35420 47124 35476
rect 47068 35028 47124 35420
rect 47068 34962 47124 34972
rect 46844 34916 46900 34926
rect 46844 34822 46900 34860
rect 46508 34804 46564 34814
rect 46396 34802 46564 34804
rect 46396 34750 46510 34802
rect 46562 34750 46564 34802
rect 46396 34748 46564 34750
rect 46396 34354 46452 34748
rect 46508 34738 46564 34748
rect 46620 34690 46676 34702
rect 46620 34638 46622 34690
rect 46674 34638 46676 34690
rect 46396 34302 46398 34354
rect 46450 34302 46452 34354
rect 46396 34290 46452 34302
rect 46508 34356 46564 34366
rect 46284 34130 46340 34142
rect 46284 34078 46286 34130
rect 46338 34078 46340 34130
rect 46284 33236 46340 34078
rect 46508 33346 46564 34300
rect 46620 33908 46676 34638
rect 47180 34692 47236 35646
rect 47404 35924 47460 35934
rect 47404 35698 47460 35868
rect 47404 35646 47406 35698
rect 47458 35646 47460 35698
rect 47404 35634 47460 35646
rect 47516 35140 47572 35150
rect 47516 34914 47572 35084
rect 47628 35028 47684 41132
rect 47852 41188 47908 41198
rect 47964 41188 48020 42702
rect 48188 42754 48244 42766
rect 48188 42702 48190 42754
rect 48242 42702 48244 42754
rect 48188 42196 48244 42702
rect 48076 41300 48132 41310
rect 48188 41300 48244 42140
rect 48412 42754 48468 42766
rect 48412 42702 48414 42754
rect 48466 42702 48468 42754
rect 48412 42084 48468 42702
rect 48412 42018 48468 42028
rect 48132 41244 48244 41300
rect 48076 41206 48132 41244
rect 47852 41186 48020 41188
rect 47852 41134 47854 41186
rect 47906 41134 48020 41186
rect 47852 41132 48020 41134
rect 47852 41076 47908 41132
rect 47852 41010 47908 41020
rect 48188 40964 48244 40974
rect 48188 40870 48244 40908
rect 48412 39620 48468 39630
rect 48412 39526 48468 39564
rect 47852 39060 47908 39070
rect 47852 38966 47908 39004
rect 48524 38668 48580 50428
rect 48860 50418 48916 50428
rect 48972 48244 49028 48254
rect 49196 48244 49252 48254
rect 48972 48150 49028 48188
rect 49084 48242 49252 48244
rect 49084 48190 49198 48242
rect 49250 48190 49252 48242
rect 49084 48188 49252 48190
rect 48860 48020 48916 48030
rect 48748 47124 48804 47134
rect 48748 46786 48804 47068
rect 48748 46734 48750 46786
rect 48802 46734 48804 46786
rect 48748 46722 48804 46734
rect 48860 46674 48916 47964
rect 48860 46622 48862 46674
rect 48914 46622 48916 46674
rect 48860 46610 48916 46622
rect 48972 47460 49028 47470
rect 48972 46564 49028 47404
rect 49084 46788 49140 48188
rect 49196 48178 49252 48188
rect 49308 46788 49364 54348
rect 49868 54292 49924 54302
rect 49868 54198 49924 54236
rect 50092 53620 50148 53630
rect 50092 53060 50148 53564
rect 50092 52946 50148 53004
rect 50092 52894 50094 52946
rect 50146 52894 50148 52946
rect 50092 52882 50148 52894
rect 50204 52276 50260 54462
rect 50652 54516 50708 54526
rect 50652 54422 50708 54460
rect 51212 54516 51268 55020
rect 51436 55298 51492 55310
rect 51436 55246 51438 55298
rect 51490 55246 51492 55298
rect 51436 54740 51492 55246
rect 52108 55188 52164 55198
rect 52668 55188 52724 55198
rect 52108 55186 52724 55188
rect 52108 55134 52110 55186
rect 52162 55134 52670 55186
rect 52722 55134 52724 55186
rect 52108 55132 52724 55134
rect 52108 55122 52164 55132
rect 52668 55122 52724 55132
rect 53004 55186 53060 56028
rect 54012 56084 54068 56094
rect 54012 55990 54068 56028
rect 53004 55134 53006 55186
rect 53058 55134 53060 55186
rect 53004 55122 53060 55134
rect 51436 54674 51492 54684
rect 51884 54740 51940 54750
rect 51884 54626 51940 54684
rect 51884 54574 51886 54626
rect 51938 54574 51940 54626
rect 51884 54562 51940 54574
rect 51660 54516 51716 54526
rect 51212 54514 51716 54516
rect 51212 54462 51214 54514
rect 51266 54462 51662 54514
rect 51714 54462 51716 54514
rect 51212 54460 51716 54462
rect 51212 54450 51268 54460
rect 51660 54450 51716 54460
rect 53228 54514 53284 54526
rect 53228 54462 53230 54514
rect 53282 54462 53284 54514
rect 50876 54404 50932 54414
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 50876 53170 50932 54348
rect 50988 54402 51044 54414
rect 50988 54350 50990 54402
rect 51042 54350 51044 54402
rect 50988 53844 51044 54350
rect 52892 54402 52948 54414
rect 52892 54350 52894 54402
rect 52946 54350 52948 54402
rect 50988 53788 51156 53844
rect 51100 53732 51156 53788
rect 51100 53666 51156 53676
rect 52780 53732 52836 53742
rect 50876 53118 50878 53170
rect 50930 53118 50932 53170
rect 50876 53106 50932 53118
rect 50988 53618 51044 53630
rect 50988 53566 50990 53618
rect 51042 53566 51044 53618
rect 50204 51492 50260 52220
rect 50316 52946 50372 52958
rect 50316 52894 50318 52946
rect 50370 52894 50372 52946
rect 50316 52052 50372 52894
rect 50428 52946 50484 52958
rect 50428 52894 50430 52946
rect 50482 52894 50484 52946
rect 50428 52164 50484 52894
rect 50428 52098 50484 52108
rect 50988 52164 51044 53566
rect 51100 53508 51156 53518
rect 51100 53506 51268 53508
rect 51100 53454 51102 53506
rect 51154 53454 51268 53506
rect 51100 53452 51268 53454
rect 51100 53442 51156 53452
rect 50988 52070 51044 52108
rect 50316 51986 50372 51996
rect 51212 52052 51268 53452
rect 51324 53506 51380 53518
rect 51324 53454 51326 53506
rect 51378 53454 51380 53506
rect 51324 52834 51380 53454
rect 51548 53060 51604 53070
rect 51604 53004 51940 53060
rect 51548 52966 51604 53004
rect 51324 52782 51326 52834
rect 51378 52782 51380 52834
rect 51324 52770 51380 52782
rect 51884 52162 51940 53004
rect 52780 52946 52836 53676
rect 52780 52894 52782 52946
rect 52834 52894 52836 52946
rect 52780 52882 52836 52894
rect 51884 52110 51886 52162
rect 51938 52110 51940 52162
rect 51884 52098 51940 52110
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 50428 51492 50484 51502
rect 50204 51490 50484 51492
rect 50204 51438 50430 51490
rect 50482 51438 50484 51490
rect 50204 51436 50484 51438
rect 50428 51426 50484 51436
rect 49420 51378 49476 51390
rect 49420 51326 49422 51378
rect 49474 51326 49476 51378
rect 49420 50484 49476 51326
rect 49644 50708 49700 50718
rect 49644 50614 49700 50652
rect 50652 50708 50708 50718
rect 50092 50596 50148 50606
rect 50092 50502 50148 50540
rect 50652 50594 50708 50652
rect 51212 50708 51268 51996
rect 51212 50642 51268 50652
rect 51996 51938 52052 51950
rect 51996 51886 51998 51938
rect 52050 51886 52052 51938
rect 51996 50708 52052 51886
rect 52892 50818 52948 54350
rect 53228 54404 53284 54462
rect 54572 54516 54628 54526
rect 54572 54422 54628 54460
rect 53228 54338 53284 54348
rect 53900 53732 53956 53742
rect 53564 53620 53620 53630
rect 53452 53618 53620 53620
rect 53452 53566 53566 53618
rect 53618 53566 53620 53618
rect 53452 53564 53620 53566
rect 53452 53058 53508 53564
rect 53564 53554 53620 53564
rect 53900 53618 53956 53676
rect 55580 53732 55636 53742
rect 55580 53638 55636 53676
rect 53900 53566 53902 53618
rect 53954 53566 53956 53618
rect 53900 53554 53956 53566
rect 57260 53618 57316 53630
rect 57260 53566 57262 53618
rect 57314 53566 57316 53618
rect 57260 53172 57316 53566
rect 57260 53106 57316 53116
rect 53452 53006 53454 53058
rect 53506 53006 53508 53058
rect 53452 52994 53508 53006
rect 55020 51492 55076 51502
rect 55020 51490 55188 51492
rect 55020 51438 55022 51490
rect 55074 51438 55188 51490
rect 55020 51436 55188 51438
rect 55020 51426 55076 51436
rect 54684 51380 54740 51390
rect 52892 50766 52894 50818
rect 52946 50766 52948 50818
rect 51996 50642 52052 50652
rect 52332 50708 52388 50718
rect 50652 50542 50654 50594
rect 50706 50542 50708 50594
rect 50652 50530 50708 50542
rect 49420 50418 49476 50428
rect 50204 50484 50260 50494
rect 50204 50390 50260 50428
rect 50764 50484 50820 50494
rect 50764 50390 50820 50428
rect 50988 50370 51044 50382
rect 50988 50318 50990 50370
rect 51042 50318 51044 50370
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 50988 49922 51044 50318
rect 50988 49870 50990 49922
rect 51042 49870 51044 49922
rect 50876 49698 50932 49710
rect 50876 49646 50878 49698
rect 50930 49646 50932 49698
rect 50876 48916 50932 49646
rect 50988 49364 51044 49870
rect 52332 49922 52388 50652
rect 52668 50708 52724 50718
rect 52668 50614 52724 50652
rect 52892 50372 52948 50766
rect 54572 51378 54740 51380
rect 54572 51326 54686 51378
rect 54738 51326 54740 51378
rect 54572 51324 54740 51326
rect 52892 50306 52948 50316
rect 53228 50708 53284 50718
rect 53676 50708 53732 50718
rect 53228 50706 53732 50708
rect 53228 50654 53230 50706
rect 53282 50654 53678 50706
rect 53730 50654 53732 50706
rect 53228 50652 53732 50654
rect 52332 49870 52334 49922
rect 52386 49870 52388 49922
rect 52332 49858 52388 49870
rect 51772 49812 51828 49822
rect 51772 49718 51828 49756
rect 53004 49812 53060 49822
rect 50988 49308 51828 49364
rect 51660 48916 51716 48926
rect 50876 48914 51716 48916
rect 50876 48862 51662 48914
rect 51714 48862 51716 48914
rect 50876 48860 51716 48862
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 49420 48356 49476 48366
rect 49420 48262 49476 48300
rect 50876 48354 50932 48860
rect 51660 48850 51716 48860
rect 51772 48914 51828 49308
rect 53004 49026 53060 49756
rect 53116 49140 53172 49150
rect 53116 49046 53172 49084
rect 53004 48974 53006 49026
rect 53058 48974 53060 49026
rect 53004 48962 53060 48974
rect 53228 49026 53284 50652
rect 53676 50642 53732 50652
rect 54572 50706 54628 51324
rect 54684 51314 54740 51324
rect 54572 50654 54574 50706
rect 54626 50654 54628 50706
rect 54572 50642 54628 50654
rect 53900 50594 53956 50606
rect 53900 50542 53902 50594
rect 53954 50542 53956 50594
rect 53900 49812 53956 50542
rect 54908 50484 54964 50494
rect 54684 50482 54964 50484
rect 54684 50430 54910 50482
rect 54962 50430 54964 50482
rect 54684 50428 54964 50430
rect 54348 50372 54404 50382
rect 53900 49718 53956 49756
rect 54236 49924 54292 49934
rect 54012 49698 54068 49710
rect 54012 49646 54014 49698
rect 54066 49646 54068 49698
rect 53900 49140 53956 49150
rect 53900 49046 53956 49084
rect 53228 48974 53230 49026
rect 53282 48974 53284 49026
rect 53228 48962 53284 48974
rect 53676 49028 53732 49038
rect 51772 48862 51774 48914
rect 51826 48862 51828 48914
rect 51772 48850 51828 48862
rect 51996 48804 52052 48814
rect 51996 48710 52052 48748
rect 52780 48804 52836 48814
rect 50876 48302 50878 48354
rect 50930 48302 50932 48354
rect 50876 48290 50932 48302
rect 50316 48242 50372 48254
rect 50316 48190 50318 48242
rect 50370 48190 50372 48242
rect 50092 48130 50148 48142
rect 50092 48078 50094 48130
rect 50146 48078 50148 48130
rect 49532 48020 49588 48030
rect 50092 48020 50148 48078
rect 49532 48018 50148 48020
rect 49532 47966 49534 48018
rect 49586 47966 50148 48018
rect 49532 47964 50148 47966
rect 49532 47954 49588 47964
rect 49532 47684 49588 47694
rect 49308 46732 49476 46788
rect 49084 46694 49140 46732
rect 49308 46564 49364 46574
rect 48972 46562 49364 46564
rect 48972 46510 49310 46562
rect 49362 46510 49364 46562
rect 48972 46508 49364 46510
rect 49308 46498 49364 46508
rect 48748 46004 48804 46014
rect 48804 45948 48916 46004
rect 48748 45938 48804 45948
rect 48748 45780 48804 45790
rect 48748 45686 48804 45724
rect 48748 45108 48804 45118
rect 48748 45014 48804 45052
rect 48860 44324 48916 45948
rect 49196 45780 49252 45790
rect 48972 45220 49028 45230
rect 48972 45126 49028 45164
rect 48860 44322 49140 44324
rect 48860 44270 48862 44322
rect 48914 44270 49140 44322
rect 48860 44268 49140 44270
rect 48860 44258 48916 44268
rect 49084 43540 49140 44268
rect 49084 43446 49140 43484
rect 48860 42532 48916 42542
rect 48860 42438 48916 42476
rect 49196 42420 49252 45724
rect 49308 45332 49364 45342
rect 49308 45218 49364 45276
rect 49308 45166 49310 45218
rect 49362 45166 49364 45218
rect 49308 45154 49364 45166
rect 49308 44436 49364 44446
rect 49420 44436 49476 46732
rect 49532 46674 49588 47628
rect 49756 47458 49812 47470
rect 49756 47406 49758 47458
rect 49810 47406 49812 47458
rect 49756 47124 49812 47406
rect 50204 47460 50260 47470
rect 50204 47366 50260 47404
rect 49756 47058 49812 47068
rect 50316 47012 50372 48190
rect 49532 46622 49534 46674
rect 49586 46622 49588 46674
rect 49532 46610 49588 46622
rect 50204 46956 50372 47012
rect 50428 48244 50484 48254
rect 50204 46674 50260 46956
rect 50316 46788 50372 46798
rect 50316 46694 50372 46732
rect 50204 46622 50206 46674
rect 50258 46622 50260 46674
rect 49980 46562 50036 46574
rect 49980 46510 49982 46562
rect 50034 46510 50036 46562
rect 49644 45780 49700 45790
rect 49980 45780 50036 46510
rect 49700 45724 50036 45780
rect 49644 45686 49700 45724
rect 49980 44996 50036 45006
rect 49980 44902 50036 44940
rect 49308 44434 49924 44436
rect 49308 44382 49310 44434
rect 49362 44382 49924 44434
rect 49308 44380 49924 44382
rect 49308 44370 49364 44380
rect 49868 43762 49924 44380
rect 49868 43710 49870 43762
rect 49922 43710 49924 43762
rect 49308 43426 49364 43438
rect 49308 43374 49310 43426
rect 49362 43374 49364 43426
rect 49308 42532 49364 43374
rect 49420 43314 49476 43326
rect 49420 43262 49422 43314
rect 49474 43262 49476 43314
rect 49420 42980 49476 43262
rect 49420 42914 49476 42924
rect 49868 42868 49924 43710
rect 50092 43764 50148 43774
rect 50204 43764 50260 46622
rect 50428 46676 50484 48188
rect 52108 48242 52164 48254
rect 52108 48190 52110 48242
rect 52162 48190 52164 48242
rect 50764 47684 50820 47694
rect 50764 47346 50820 47628
rect 52108 47460 52164 48190
rect 52108 47348 52164 47404
rect 50764 47294 50766 47346
rect 50818 47294 50820 47346
rect 50764 47282 50820 47294
rect 51884 47292 52164 47348
rect 52444 48244 52500 48254
rect 51772 47236 51828 47246
rect 51772 47142 51828 47180
rect 50988 47124 51044 47134
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 50988 46898 51044 47068
rect 50988 46846 50990 46898
rect 51042 46846 51044 46898
rect 50988 46834 51044 46846
rect 50540 46676 50596 46686
rect 50428 46674 50596 46676
rect 50428 46622 50542 46674
rect 50594 46622 50596 46674
rect 50428 46620 50596 46622
rect 50540 46610 50596 46620
rect 51772 46676 51828 46686
rect 51884 46676 51940 47292
rect 52220 47236 52276 47246
rect 52444 47236 52500 48188
rect 52668 48242 52724 48254
rect 52668 48190 52670 48242
rect 52722 48190 52724 48242
rect 52276 47180 52500 47236
rect 52556 48130 52612 48142
rect 52556 48078 52558 48130
rect 52610 48078 52612 48130
rect 51772 46674 51940 46676
rect 51772 46622 51774 46674
rect 51826 46622 51940 46674
rect 51772 46620 51940 46622
rect 51996 47124 52052 47134
rect 51996 46674 52052 47068
rect 51996 46622 51998 46674
rect 52050 46622 52052 46674
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 50316 45220 50372 45230
rect 50316 45106 50372 45164
rect 50316 45054 50318 45106
rect 50370 45054 50372 45106
rect 50316 45042 50372 45054
rect 50988 45106 51044 45118
rect 50988 45054 50990 45106
rect 51042 45054 51044 45106
rect 50764 44996 50820 45006
rect 50652 44436 50708 44446
rect 50764 44436 50820 44940
rect 50876 44436 50932 44446
rect 50764 44434 50932 44436
rect 50764 44382 50878 44434
rect 50930 44382 50932 44434
rect 50764 44380 50932 44382
rect 50652 44322 50708 44380
rect 50876 44370 50932 44380
rect 50988 44436 51044 45054
rect 50988 44370 51044 44380
rect 51212 44882 51268 44894
rect 51212 44830 51214 44882
rect 51266 44830 51268 44882
rect 50652 44270 50654 44322
rect 50706 44270 50708 44322
rect 50652 44258 50708 44270
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 50148 43708 50260 43764
rect 50092 43698 50148 43708
rect 51212 43652 51268 44830
rect 51324 44436 51380 44446
rect 51772 44436 51828 46620
rect 51996 46610 52052 46622
rect 52220 46674 52276 47180
rect 52220 46622 52222 46674
rect 52274 46622 52276 46674
rect 52220 46610 52276 46622
rect 52332 46676 52388 46686
rect 52556 46676 52612 48078
rect 52668 48020 52724 48190
rect 52668 47124 52724 47964
rect 52668 47058 52724 47068
rect 52780 46786 52836 48748
rect 53228 48354 53284 48366
rect 53228 48302 53230 48354
rect 53282 48302 53284 48354
rect 53228 48244 53284 48302
rect 53228 48178 53284 48188
rect 53116 48130 53172 48142
rect 53116 48078 53118 48130
rect 53170 48078 53172 48130
rect 53004 48020 53060 48030
rect 53004 47926 53060 47964
rect 52892 47570 52948 47582
rect 52892 47518 52894 47570
rect 52946 47518 52948 47570
rect 52892 47460 52948 47518
rect 52892 47394 52948 47404
rect 53116 47458 53172 48078
rect 53676 47570 53732 48972
rect 53676 47518 53678 47570
rect 53730 47518 53732 47570
rect 53676 47506 53732 47518
rect 53116 47406 53118 47458
rect 53170 47406 53172 47458
rect 53116 47394 53172 47406
rect 52780 46734 52782 46786
rect 52834 46734 52836 46786
rect 52780 46722 52836 46734
rect 53676 46898 53732 46910
rect 53676 46846 53678 46898
rect 53730 46846 53732 46898
rect 52668 46676 52724 46686
rect 52556 46674 52724 46676
rect 52556 46622 52670 46674
rect 52722 46622 52724 46674
rect 52556 46620 52724 46622
rect 52332 46582 52388 46620
rect 52668 46610 52724 46620
rect 53564 46676 53620 46686
rect 53564 46582 53620 46620
rect 53564 45220 53620 45230
rect 53676 45220 53732 46846
rect 53564 45218 53732 45220
rect 53564 45166 53566 45218
rect 53618 45166 53732 45218
rect 53564 45164 53732 45166
rect 53564 45154 53620 45164
rect 51324 44434 51828 44436
rect 51324 44382 51326 44434
rect 51378 44382 51828 44434
rect 51324 44380 51828 44382
rect 53676 44434 53732 45164
rect 53676 44382 53678 44434
rect 53730 44382 53732 44434
rect 51324 44370 51380 44380
rect 53676 44370 53732 44382
rect 53788 45332 53844 45342
rect 54012 45332 54068 49646
rect 54236 49028 54292 49868
rect 54348 49810 54404 50316
rect 54348 49758 54350 49810
rect 54402 49758 54404 49810
rect 54348 49746 54404 49758
rect 54236 48934 54292 48972
rect 54684 49026 54740 50428
rect 54908 50418 54964 50428
rect 54908 49924 54964 49934
rect 54908 49830 54964 49868
rect 55132 49140 55188 51436
rect 57932 50706 57988 50718
rect 57932 50654 57934 50706
rect 57986 50654 57988 50706
rect 55580 50596 55636 50606
rect 55244 50594 55636 50596
rect 55244 50542 55582 50594
rect 55634 50542 55636 50594
rect 55244 50540 55636 50542
rect 55244 50482 55300 50540
rect 55580 50530 55636 50540
rect 55244 50430 55246 50482
rect 55298 50430 55300 50482
rect 55244 50418 55300 50430
rect 57820 50372 57876 50382
rect 55132 49084 55300 49140
rect 54684 48974 54686 49026
rect 54738 48974 54740 49026
rect 54684 48962 54740 48974
rect 55244 49028 55300 49084
rect 57820 49138 57876 50316
rect 57932 49812 57988 50654
rect 57932 49746 57988 49756
rect 57820 49086 57822 49138
rect 57874 49086 57876 49138
rect 57820 49074 57876 49086
rect 55580 49028 55636 49038
rect 55244 49026 55636 49028
rect 55244 48974 55582 49026
rect 55634 48974 55636 49026
rect 55244 48972 55636 48974
rect 55580 48962 55636 48972
rect 58156 47234 58212 47246
rect 58156 47182 58158 47234
rect 58210 47182 58212 47234
rect 58156 47124 58212 47182
rect 58156 47058 58212 47068
rect 53788 45330 54068 45332
rect 53788 45278 53790 45330
rect 53842 45278 54068 45330
rect 53788 45276 54068 45278
rect 53116 44324 53172 44334
rect 51212 43586 51268 43596
rect 51436 43650 51492 43662
rect 51436 43598 51438 43650
rect 51490 43598 51492 43650
rect 51324 43538 51380 43550
rect 51324 43486 51326 43538
rect 51378 43486 51380 43538
rect 49420 42756 49476 42766
rect 49420 42662 49476 42700
rect 49308 42476 49476 42532
rect 48972 42364 49252 42420
rect 48748 41970 48804 41982
rect 48748 41918 48750 41970
rect 48802 41918 48804 41970
rect 48636 41188 48692 41198
rect 48636 41094 48692 41132
rect 48748 41076 48804 41918
rect 48972 41972 49028 42364
rect 49084 42196 49140 42206
rect 49084 42102 49140 42140
rect 49308 42084 49364 42094
rect 49308 41990 49364 42028
rect 49196 41972 49252 41982
rect 49028 41916 49140 41972
rect 48972 41906 49028 41916
rect 49084 41300 49140 41916
rect 49420 41972 49476 42476
rect 49756 41972 49812 41982
rect 49420 41970 49812 41972
rect 49420 41918 49758 41970
rect 49810 41918 49812 41970
rect 49420 41916 49812 41918
rect 49196 41878 49252 41916
rect 49756 41906 49812 41916
rect 49868 41748 49924 42812
rect 49980 42980 50036 42990
rect 49980 42642 50036 42924
rect 51212 42868 51268 42878
rect 51212 42774 51268 42812
rect 49980 42590 49982 42642
rect 50034 42590 50036 42642
rect 49980 42578 50036 42590
rect 50092 42756 50148 42766
rect 50092 41970 50148 42700
rect 50876 42532 50932 42542
rect 50092 41918 50094 41970
rect 50146 41918 50148 41970
rect 50092 41906 50148 41918
rect 50428 42530 50932 42532
rect 50428 42478 50878 42530
rect 50930 42478 50932 42530
rect 50428 42476 50932 42478
rect 49644 41692 49924 41748
rect 49140 41244 49252 41300
rect 49084 41206 49140 41244
rect 48748 41010 48804 41020
rect 48860 40404 48916 40414
rect 48748 40402 48916 40404
rect 48748 40350 48862 40402
rect 48914 40350 48916 40402
rect 48748 40348 48916 40350
rect 48636 39618 48692 39630
rect 48636 39566 48638 39618
rect 48690 39566 48692 39618
rect 48636 39396 48692 39566
rect 48636 39330 48692 39340
rect 47628 34962 47684 34972
rect 47740 38612 48580 38668
rect 48748 38724 48804 40348
rect 48860 40338 48916 40348
rect 49084 39844 49140 39854
rect 48972 39508 49028 39518
rect 48972 39414 49028 39452
rect 48972 39060 49028 39070
rect 48972 38834 49028 39004
rect 48972 38782 48974 38834
rect 49026 38782 49028 38834
rect 48972 38770 49028 38782
rect 49084 38836 49140 39788
rect 49196 39730 49252 41244
rect 49420 40516 49476 40526
rect 49420 40422 49476 40460
rect 49196 39678 49198 39730
rect 49250 39678 49252 39730
rect 49196 39666 49252 39678
rect 49308 40402 49364 40414
rect 49308 40350 49310 40402
rect 49362 40350 49364 40402
rect 49308 39060 49364 40350
rect 49532 40402 49588 40414
rect 49532 40350 49534 40402
rect 49586 40350 49588 40402
rect 49532 39844 49588 40350
rect 49532 39778 49588 39788
rect 49644 39508 49700 41692
rect 49980 41300 50036 41310
rect 49980 40626 50036 41244
rect 49980 40574 49982 40626
rect 50034 40574 50036 40626
rect 49980 40562 50036 40574
rect 49756 39842 49812 39854
rect 49756 39790 49758 39842
rect 49810 39790 49812 39842
rect 49756 39620 49812 39790
rect 49756 39554 49812 39564
rect 49868 39730 49924 39742
rect 49868 39678 49870 39730
rect 49922 39678 49924 39730
rect 49644 39414 49700 39452
rect 49868 39396 49924 39678
rect 49868 39330 49924 39340
rect 50092 39508 50148 39518
rect 49308 38994 49364 39004
rect 49644 39060 49700 39070
rect 49644 38966 49700 39004
rect 50092 39058 50148 39452
rect 50092 39006 50094 39058
rect 50146 39006 50148 39058
rect 50092 38948 50148 39006
rect 50092 38882 50148 38892
rect 49196 38836 49252 38846
rect 49084 38834 49252 38836
rect 49084 38782 49198 38834
rect 49250 38782 49252 38834
rect 49084 38780 49252 38782
rect 49196 38770 49252 38780
rect 48748 38658 48804 38668
rect 47516 34862 47518 34914
rect 47570 34862 47572 34914
rect 47516 34850 47572 34862
rect 47180 34636 47684 34692
rect 46844 34356 46900 34366
rect 46844 34242 46900 34300
rect 46844 34190 46846 34242
rect 46898 34190 46900 34242
rect 46844 34178 46900 34190
rect 46956 34242 47012 34254
rect 46956 34190 46958 34242
rect 47010 34190 47012 34242
rect 46956 34132 47012 34190
rect 47628 34242 47684 34636
rect 47628 34190 47630 34242
rect 47682 34190 47684 34242
rect 47628 34178 47684 34190
rect 46956 34076 47124 34132
rect 46956 33908 47012 33918
rect 46620 33906 47012 33908
rect 46620 33854 46958 33906
rect 47010 33854 47012 33906
rect 46620 33852 47012 33854
rect 46956 33842 47012 33852
rect 46508 33294 46510 33346
rect 46562 33294 46564 33346
rect 46508 33282 46564 33294
rect 46284 33170 46340 33180
rect 47068 33236 47124 34076
rect 47516 33460 47572 33470
rect 47180 33348 47236 33358
rect 47516 33348 47572 33404
rect 47180 33254 47236 33292
rect 47292 33346 47572 33348
rect 47292 33294 47518 33346
rect 47570 33294 47572 33346
rect 47292 33292 47572 33294
rect 47068 33170 47124 33180
rect 46956 32676 47012 32686
rect 46956 32582 47012 32620
rect 47180 32564 47236 32574
rect 47292 32564 47348 33292
rect 47516 33282 47572 33292
rect 47628 33122 47684 33134
rect 47628 33070 47630 33122
rect 47682 33070 47684 33122
rect 47516 32788 47572 32798
rect 47516 32694 47572 32732
rect 47628 32676 47684 33070
rect 47628 32610 47684 32620
rect 47180 32562 47348 32564
rect 47180 32510 47182 32562
rect 47234 32510 47348 32562
rect 47180 32508 47348 32510
rect 47180 32498 47236 32508
rect 46172 31838 46174 31890
rect 46226 31838 46228 31890
rect 46172 31220 46228 31838
rect 46172 31218 46788 31220
rect 46172 31166 46174 31218
rect 46226 31166 46788 31218
rect 46172 31164 46788 31166
rect 46172 31154 46228 31164
rect 46508 30996 46564 31006
rect 45948 30994 46564 30996
rect 45948 30942 46510 30994
rect 46562 30942 46564 30994
rect 45948 30940 46564 30942
rect 45948 30210 46004 30940
rect 45948 30158 45950 30210
rect 46002 30158 46004 30210
rect 45948 30146 46004 30158
rect 45836 30046 45838 30098
rect 45890 30046 45892 30098
rect 45836 30034 45892 30046
rect 43932 29986 43988 29998
rect 43932 29934 43934 29986
rect 43986 29934 43988 29986
rect 43932 29428 43988 29934
rect 46396 29650 46452 30940
rect 46508 30930 46564 30940
rect 46732 30994 46788 31164
rect 47292 31108 47348 31118
rect 47740 31108 47796 38612
rect 50428 37492 50484 42476
rect 50876 42466 50932 42476
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 51212 41972 51268 41982
rect 51324 41972 51380 43486
rect 51436 42532 51492 43598
rect 51772 43652 51828 43662
rect 51660 43540 51716 43550
rect 51660 43446 51716 43484
rect 51772 42756 51828 43596
rect 52220 43652 52276 43662
rect 52220 43538 52276 43596
rect 53116 43650 53172 44268
rect 53788 44322 53844 45276
rect 55916 45218 55972 45230
rect 55916 45166 55918 45218
rect 55970 45166 55972 45218
rect 54572 45108 54628 45118
rect 54460 45106 54628 45108
rect 54460 45054 54574 45106
rect 54626 45054 54628 45106
rect 54460 45052 54628 45054
rect 53900 44996 53956 45006
rect 54348 44996 54404 45006
rect 53900 44994 54404 44996
rect 53900 44942 53902 44994
rect 53954 44942 54350 44994
rect 54402 44942 54404 44994
rect 53900 44940 54404 44942
rect 53900 44930 53956 44940
rect 53788 44270 53790 44322
rect 53842 44270 53844 44322
rect 53788 44258 53844 44270
rect 54124 43762 54180 44940
rect 54348 44930 54404 44940
rect 54124 43710 54126 43762
rect 54178 43710 54180 43762
rect 54124 43698 54180 43710
rect 53900 43652 53956 43662
rect 53116 43598 53118 43650
rect 53170 43598 53172 43650
rect 53116 43586 53172 43598
rect 53676 43596 53900 43652
rect 52220 43486 52222 43538
rect 52274 43486 52276 43538
rect 52220 43474 52276 43486
rect 52332 43540 52388 43550
rect 52332 43428 52388 43484
rect 52892 43540 52948 43550
rect 52332 43426 52836 43428
rect 52332 43374 52334 43426
rect 52386 43374 52836 43426
rect 52332 43372 52836 43374
rect 52332 43362 52388 43372
rect 52780 42866 52836 43372
rect 52780 42814 52782 42866
rect 52834 42814 52836 42866
rect 52780 42802 52836 42814
rect 51548 42532 51604 42542
rect 51436 42476 51548 42532
rect 51548 42194 51604 42476
rect 51548 42142 51550 42194
rect 51602 42142 51604 42194
rect 51548 42130 51604 42142
rect 51772 42194 51828 42700
rect 51772 42142 51774 42194
rect 51826 42142 51828 42194
rect 51772 42130 51828 42142
rect 51884 42196 51940 42206
rect 51268 41916 51380 41972
rect 51436 41972 51492 41982
rect 51212 41878 51268 41916
rect 50652 41860 50708 41870
rect 50652 41858 50932 41860
rect 50652 41806 50654 41858
rect 50706 41806 50932 41858
rect 50652 41804 50932 41806
rect 50652 41794 50708 41804
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 50540 40516 50596 40526
rect 50540 40422 50596 40460
rect 50764 40402 50820 40414
rect 50764 40350 50766 40402
rect 50818 40350 50820 40402
rect 50764 39956 50820 40350
rect 50764 39890 50820 39900
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 50540 38948 50596 38958
rect 50540 38854 50596 38892
rect 50876 38052 50932 41804
rect 51324 41074 51380 41086
rect 51324 41022 51326 41074
rect 51378 41022 51380 41074
rect 50988 40964 51044 40974
rect 51324 40964 51380 41022
rect 51044 40908 51380 40964
rect 50988 40626 51044 40908
rect 50988 40574 50990 40626
rect 51042 40574 51044 40626
rect 50988 40562 51044 40574
rect 51324 40402 51380 40908
rect 51324 40350 51326 40402
rect 51378 40350 51380 40402
rect 51324 40338 51380 40350
rect 51100 40180 51156 40190
rect 51436 40180 51492 41916
rect 51884 41970 51940 42140
rect 52556 42196 52612 42206
rect 52556 42102 52612 42140
rect 51884 41918 51886 41970
rect 51938 41918 51940 41970
rect 51884 41906 51940 41918
rect 52444 41972 52500 41982
rect 52444 41878 52500 41916
rect 52780 41970 52836 41982
rect 52780 41918 52782 41970
rect 52834 41918 52836 41970
rect 52668 41188 52724 41198
rect 52108 41186 52724 41188
rect 52108 41134 52670 41186
rect 52722 41134 52724 41186
rect 52108 41132 52724 41134
rect 51100 40178 51492 40180
rect 51100 40126 51102 40178
rect 51154 40126 51492 40178
rect 51100 40124 51492 40126
rect 51548 41074 51604 41086
rect 51548 41022 51550 41074
rect 51602 41022 51604 41074
rect 51548 40402 51604 41022
rect 51772 41076 51828 41086
rect 51772 40982 51828 41020
rect 51884 41074 51940 41086
rect 51884 41022 51886 41074
rect 51938 41022 51940 41074
rect 51660 40516 51716 40526
rect 51884 40516 51940 41022
rect 52108 40626 52164 41132
rect 52668 41122 52724 41132
rect 52780 40740 52836 41918
rect 52892 41298 52948 43484
rect 53452 43538 53508 43550
rect 53452 43486 53454 43538
rect 53506 43486 53508 43538
rect 53004 42756 53060 42766
rect 53004 42662 53060 42700
rect 53452 42196 53508 43486
rect 53676 42866 53732 43596
rect 53900 43558 53956 43596
rect 54460 43652 54516 45052
rect 54572 45042 54628 45052
rect 55244 45108 55300 45118
rect 55580 45108 55636 45118
rect 55244 45106 55636 45108
rect 55244 45054 55246 45106
rect 55298 45054 55582 45106
rect 55634 45054 55636 45106
rect 55244 45052 55636 45054
rect 55244 45042 55300 45052
rect 55580 45042 55636 45052
rect 54684 44434 54740 44446
rect 54684 44382 54686 44434
rect 54738 44382 54740 44434
rect 54572 44324 54628 44334
rect 54572 44230 54628 44268
rect 54460 43586 54516 43596
rect 54012 43428 54068 43438
rect 54572 43428 54628 43438
rect 54012 43426 54628 43428
rect 54012 43374 54014 43426
rect 54066 43374 54574 43426
rect 54626 43374 54628 43426
rect 54012 43372 54628 43374
rect 54012 43362 54068 43372
rect 54572 43362 54628 43372
rect 53676 42814 53678 42866
rect 53730 42814 53732 42866
rect 53676 42802 53732 42814
rect 53452 42130 53508 42140
rect 52892 41246 52894 41298
rect 52946 41246 52948 41298
rect 52892 41234 52948 41246
rect 54572 41188 54628 41198
rect 54684 41188 54740 44382
rect 55916 44322 55972 45166
rect 57932 44436 57988 44446
rect 57932 44342 57988 44380
rect 55916 44270 55918 44322
rect 55970 44270 55972 44322
rect 55916 44258 55972 44270
rect 54908 44210 54964 44222
rect 54908 44158 54910 44210
rect 54962 44158 54964 44210
rect 54908 43708 54964 44158
rect 54796 43652 54964 43708
rect 56588 43652 56644 43662
rect 54796 43540 54852 43652
rect 56028 43650 56644 43652
rect 56028 43598 56590 43650
rect 56642 43598 56644 43650
rect 56028 43596 56644 43598
rect 54796 43446 54852 43484
rect 55468 43540 55524 43550
rect 55468 43446 55524 43484
rect 56028 42754 56084 43596
rect 56588 43586 56644 43596
rect 56812 43540 56868 43550
rect 56812 43446 56868 43484
rect 57932 43092 57988 43102
rect 57932 42978 57988 43036
rect 57932 42926 57934 42978
rect 57986 42926 57988 42978
rect 57932 42914 57988 42926
rect 56028 42702 56030 42754
rect 56082 42702 56084 42754
rect 56028 42690 56084 42702
rect 57932 41298 57988 41310
rect 57932 41246 57934 41298
rect 57986 41246 57988 41298
rect 54572 41186 54740 41188
rect 54572 41134 54574 41186
rect 54626 41134 54740 41186
rect 54572 41132 54740 41134
rect 56028 41186 56084 41198
rect 56028 41134 56030 41186
rect 56082 41134 56084 41186
rect 53004 41076 53060 41086
rect 53340 41076 53396 41086
rect 53060 41074 53396 41076
rect 53060 41022 53342 41074
rect 53394 41022 53396 41074
rect 53060 41020 53396 41022
rect 53004 40982 53060 41020
rect 53340 41010 53396 41020
rect 54348 41076 54404 41086
rect 54348 40982 54404 41020
rect 54460 41074 54516 41086
rect 54460 41022 54462 41074
rect 54514 41022 54516 41074
rect 53452 40962 53508 40974
rect 53452 40910 53454 40962
rect 53506 40910 53508 40962
rect 52780 40684 53396 40740
rect 52108 40574 52110 40626
rect 52162 40574 52164 40626
rect 52108 40562 52164 40574
rect 51716 40460 51940 40516
rect 53340 40514 53396 40684
rect 53452 40626 53508 40910
rect 53452 40574 53454 40626
rect 53506 40574 53508 40626
rect 53452 40562 53508 40574
rect 53676 40628 53732 40638
rect 53676 40534 53732 40572
rect 54460 40628 54516 41022
rect 53340 40462 53342 40514
rect 53394 40462 53396 40514
rect 51660 40422 51716 40460
rect 53340 40450 53396 40462
rect 54460 40514 54516 40572
rect 54460 40462 54462 40514
rect 54514 40462 54516 40514
rect 54460 40450 54516 40462
rect 51548 40350 51550 40402
rect 51602 40350 51604 40402
rect 51100 40114 51156 40124
rect 51100 39956 51156 39966
rect 51548 39956 51604 40350
rect 54572 40402 54628 41132
rect 55132 41076 55188 41086
rect 54572 40350 54574 40402
rect 54626 40350 54628 40402
rect 54572 40338 54628 40350
rect 55020 40962 55076 40974
rect 55020 40910 55022 40962
rect 55074 40910 55076 40962
rect 55020 40292 55076 40910
rect 55020 40226 55076 40236
rect 55132 40402 55188 41020
rect 55132 40350 55134 40402
rect 55186 40350 55188 40402
rect 51156 39900 51604 39956
rect 51100 39618 51156 39900
rect 54124 39842 54180 39854
rect 54124 39790 54126 39842
rect 54178 39790 54180 39842
rect 54124 39732 54180 39790
rect 54124 39676 54516 39732
rect 51100 39566 51102 39618
rect 51154 39566 51156 39618
rect 50988 39508 51044 39518
rect 50988 39414 51044 39452
rect 51100 39060 51156 39566
rect 51100 38994 51156 39004
rect 53228 39508 53284 39518
rect 53228 39060 53284 39452
rect 54236 39506 54292 39518
rect 54236 39454 54238 39506
rect 54290 39454 54292 39506
rect 54124 39396 54180 39406
rect 53228 38966 53284 39004
rect 53900 39394 54180 39396
rect 53900 39342 54126 39394
rect 54178 39342 54180 39394
rect 53900 39340 54180 39342
rect 51884 38836 51940 38846
rect 51436 38162 51492 38174
rect 51436 38110 51438 38162
rect 51490 38110 51492 38162
rect 51212 38052 51268 38062
rect 50876 38050 51268 38052
rect 50876 37998 51214 38050
rect 51266 37998 51268 38050
rect 50876 37996 51268 37998
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 50540 37492 50596 37502
rect 50428 37490 50596 37492
rect 50428 37438 50542 37490
rect 50594 37438 50596 37490
rect 50428 37436 50596 37438
rect 49756 37380 49812 37390
rect 49756 37286 49812 37324
rect 50092 37268 50148 37278
rect 49868 37156 49924 37166
rect 49868 37062 49924 37100
rect 49308 36594 49364 36606
rect 49308 36542 49310 36594
rect 49362 36542 49364 36594
rect 48524 36484 48580 36494
rect 47964 36482 48580 36484
rect 47964 36430 48526 36482
rect 48578 36430 48580 36482
rect 47964 36428 48580 36430
rect 47852 35924 47908 35934
rect 47852 34354 47908 35868
rect 47852 34302 47854 34354
rect 47906 34302 47908 34354
rect 47852 34290 47908 34302
rect 47964 34018 48020 36428
rect 48524 36418 48580 36428
rect 49196 36370 49252 36382
rect 49196 36318 49198 36370
rect 49250 36318 49252 36370
rect 48076 35812 48132 35822
rect 48076 35718 48132 35756
rect 49084 35700 49140 35710
rect 49196 35700 49252 36318
rect 49140 35644 49252 35700
rect 49084 35606 49140 35644
rect 48860 35476 48916 35486
rect 48860 35138 48916 35420
rect 48860 35086 48862 35138
rect 48914 35086 48916 35138
rect 48860 35074 48916 35086
rect 49308 35140 49364 36542
rect 49532 36482 49588 36494
rect 49532 36430 49534 36482
rect 49586 36430 49588 36482
rect 49532 35812 49588 36430
rect 49532 35698 49588 35756
rect 49756 35812 49812 35822
rect 50092 35812 50148 37212
rect 50540 37268 50596 37436
rect 50652 37492 50708 37502
rect 50652 37398 50708 37436
rect 50540 37202 50596 37212
rect 50764 37268 50820 37278
rect 51100 37268 51156 37278
rect 50764 37266 51156 37268
rect 50764 37214 50766 37266
rect 50818 37214 51102 37266
rect 51154 37214 51156 37266
rect 50764 37212 51156 37214
rect 50764 37202 50820 37212
rect 50988 36706 51044 37212
rect 51100 37202 51156 37212
rect 50988 36654 50990 36706
rect 51042 36654 51044 36706
rect 50988 36642 51044 36654
rect 51212 36482 51268 37996
rect 51436 37156 51492 38110
rect 51884 38162 51940 38780
rect 53116 38836 53172 38846
rect 53116 38742 53172 38780
rect 53452 38836 53508 38846
rect 53452 38834 53732 38836
rect 53452 38782 53454 38834
rect 53506 38782 53732 38834
rect 53452 38780 53732 38782
rect 53452 38770 53508 38780
rect 53228 38276 53284 38286
rect 53228 38274 53396 38276
rect 53228 38222 53230 38274
rect 53282 38222 53396 38274
rect 53228 38220 53396 38222
rect 53228 38210 53284 38220
rect 51884 38110 51886 38162
rect 51938 38110 51940 38162
rect 51884 38098 51940 38110
rect 51660 37380 51716 37390
rect 51660 37286 51716 37324
rect 52892 37268 52948 37278
rect 52892 37174 52948 37212
rect 51436 36594 51492 37100
rect 51436 36542 51438 36594
rect 51490 36542 51492 36594
rect 51436 36530 51492 36542
rect 53004 37154 53060 37166
rect 53004 37102 53006 37154
rect 53058 37102 53060 37154
rect 51212 36430 51214 36482
rect 51266 36430 51268 36482
rect 51212 36418 51268 36430
rect 53004 36372 53060 37102
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 49756 35810 50148 35812
rect 49756 35758 49758 35810
rect 49810 35758 50148 35810
rect 49756 35756 50148 35758
rect 49756 35746 49812 35756
rect 52556 35700 52612 35710
rect 49532 35646 49534 35698
rect 49586 35646 49588 35698
rect 49532 35634 49588 35646
rect 52444 35698 52612 35700
rect 52444 35646 52558 35698
rect 52610 35646 52612 35698
rect 52444 35644 52612 35646
rect 49308 35074 49364 35084
rect 50428 35140 50484 35150
rect 48076 35028 48132 35038
rect 48076 34914 48132 34972
rect 50316 35028 50372 35038
rect 50316 34934 50372 34972
rect 48076 34862 48078 34914
rect 48130 34862 48132 34914
rect 48076 34850 48132 34862
rect 48748 34916 48804 34926
rect 48748 34822 48804 34860
rect 49196 34914 49252 34926
rect 49196 34862 49198 34914
rect 49250 34862 49252 34914
rect 49196 34692 49252 34862
rect 49420 34916 49476 34926
rect 49756 34916 49812 34926
rect 49420 34914 49812 34916
rect 49420 34862 49422 34914
rect 49474 34862 49758 34914
rect 49810 34862 49812 34914
rect 49420 34860 49812 34862
rect 49420 34850 49476 34860
rect 49756 34850 49812 34860
rect 49196 34626 49252 34636
rect 49868 34802 49924 34814
rect 49868 34750 49870 34802
rect 49922 34750 49924 34802
rect 49868 34354 49924 34750
rect 49868 34302 49870 34354
rect 49922 34302 49924 34354
rect 49868 34290 49924 34302
rect 50428 34244 50484 35084
rect 51996 34804 52052 34814
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 50876 34356 50932 34366
rect 50876 34262 50932 34300
rect 51436 34356 51492 34366
rect 50652 34244 50708 34254
rect 50428 34188 50652 34244
rect 50652 34150 50708 34188
rect 49644 34132 49700 34142
rect 47964 33966 47966 34018
rect 48018 33966 48020 34018
rect 47964 33954 48020 33966
rect 49308 34130 49700 34132
rect 49308 34078 49646 34130
rect 49698 34078 49700 34130
rect 49308 34076 49700 34078
rect 49308 33570 49364 34076
rect 49644 34066 49700 34076
rect 50092 34132 50148 34142
rect 50092 34038 50148 34076
rect 50204 34130 50260 34142
rect 50204 34078 50206 34130
rect 50258 34078 50260 34130
rect 50204 33572 50260 34078
rect 50764 34132 50820 34142
rect 50764 34038 50820 34076
rect 49308 33518 49310 33570
rect 49362 33518 49364 33570
rect 49308 33506 49364 33518
rect 49980 33516 50260 33572
rect 49980 33458 50036 33516
rect 49980 33406 49982 33458
rect 50034 33406 50036 33458
rect 49980 33394 50036 33406
rect 48636 33348 48692 33358
rect 48636 33254 48692 33292
rect 49532 33348 49588 33358
rect 48188 33236 48244 33246
rect 47852 33124 47908 33134
rect 47852 33122 48020 33124
rect 47852 33070 47854 33122
rect 47906 33070 48020 33122
rect 47852 33068 48020 33070
rect 47852 33058 47908 33068
rect 47964 32674 48020 33068
rect 48076 32788 48132 32798
rect 48076 32694 48132 32732
rect 47964 32622 47966 32674
rect 48018 32622 48020 32674
rect 47964 32610 48020 32622
rect 48188 32004 48244 33180
rect 48524 33236 48580 33246
rect 48524 33142 48580 33180
rect 48188 31938 48244 31948
rect 48300 33122 48356 33134
rect 48300 33070 48302 33122
rect 48354 33070 48356 33122
rect 48300 32562 48356 33070
rect 48300 32510 48302 32562
rect 48354 32510 48356 32562
rect 48300 31892 48356 32510
rect 48972 33122 49028 33134
rect 48972 33070 48974 33122
rect 49026 33070 49028 33122
rect 48860 32004 48916 32014
rect 48972 32004 49028 33070
rect 49196 33122 49252 33134
rect 49196 33070 49198 33122
rect 49250 33070 49252 33122
rect 49196 32788 49252 33070
rect 49196 32722 49252 32732
rect 49532 32564 49588 33292
rect 50204 33348 50260 33516
rect 51436 33570 51492 34300
rect 51996 34354 52052 34748
rect 51996 34302 51998 34354
rect 52050 34302 52052 34354
rect 51996 34290 52052 34302
rect 52444 34244 52500 35644
rect 52556 35634 52612 35644
rect 52780 35700 52836 35710
rect 52780 35698 52948 35700
rect 52780 35646 52782 35698
rect 52834 35646 52948 35698
rect 52780 35644 52948 35646
rect 52780 35634 52836 35644
rect 52668 35586 52724 35598
rect 52668 35534 52670 35586
rect 52722 35534 52724 35586
rect 52668 35140 52724 35534
rect 52556 35084 52724 35140
rect 52780 35252 52836 35262
rect 52556 34468 52612 35084
rect 52780 35028 52836 35196
rect 52668 34972 52836 35028
rect 52668 34914 52724 34972
rect 52668 34862 52670 34914
rect 52722 34862 52724 34914
rect 52668 34850 52724 34862
rect 52892 34916 52948 35644
rect 53004 35698 53060 36316
rect 53004 35646 53006 35698
rect 53058 35646 53060 35698
rect 53004 35634 53060 35646
rect 53228 35700 53284 35710
rect 53228 35606 53284 35644
rect 53340 35700 53396 38220
rect 53564 38162 53620 38174
rect 53564 38110 53566 38162
rect 53618 38110 53620 38162
rect 53452 38052 53508 38062
rect 53452 37958 53508 37996
rect 53564 36482 53620 38110
rect 53676 37380 53732 38780
rect 53900 37492 53956 39340
rect 54124 39330 54180 39340
rect 54124 39060 54180 39070
rect 53676 37324 53844 37380
rect 53564 36430 53566 36482
rect 53618 36430 53620 36482
rect 53564 36418 53620 36430
rect 53788 36370 53844 37324
rect 53900 36482 53956 37436
rect 54012 38836 54068 38846
rect 54012 38722 54068 38780
rect 54124 38834 54180 39004
rect 54124 38782 54126 38834
rect 54178 38782 54180 38834
rect 54124 38770 54180 38782
rect 54012 38670 54014 38722
rect 54066 38670 54068 38722
rect 54012 37380 54068 38670
rect 54012 37324 54180 37380
rect 54124 37266 54180 37324
rect 54124 37214 54126 37266
rect 54178 37214 54180 37266
rect 54124 37202 54180 37214
rect 54236 36706 54292 39454
rect 54348 38050 54404 38062
rect 54348 37998 54350 38050
rect 54402 37998 54404 38050
rect 54348 37490 54404 37998
rect 54460 38052 54516 39676
rect 54572 39060 54628 39070
rect 54628 39004 54740 39060
rect 54572 38994 54628 39004
rect 54572 38052 54628 38062
rect 54460 38050 54628 38052
rect 54460 37998 54574 38050
rect 54626 37998 54628 38050
rect 54460 37996 54628 37998
rect 54572 37986 54628 37996
rect 54348 37438 54350 37490
rect 54402 37438 54404 37490
rect 54348 37426 54404 37438
rect 54572 37380 54628 37390
rect 54684 37380 54740 39004
rect 54796 38948 54852 38958
rect 55132 38948 55188 40350
rect 54796 38946 55188 38948
rect 54796 38894 54798 38946
rect 54850 38894 55188 38946
rect 54796 38892 55188 38894
rect 55244 40626 55300 40638
rect 55244 40574 55246 40626
rect 55298 40574 55300 40626
rect 55244 40404 55300 40574
rect 56028 40516 56084 41134
rect 56588 40516 56644 40526
rect 56028 40514 56644 40516
rect 56028 40462 56590 40514
rect 56642 40462 56644 40514
rect 56028 40460 56644 40462
rect 56588 40450 56644 40460
rect 54796 38882 54852 38892
rect 55244 38724 55300 40348
rect 56924 40404 56980 40414
rect 56924 40310 56980 40348
rect 57932 40404 57988 41246
rect 57932 40338 57988 40348
rect 56812 40292 56868 40302
rect 56812 40198 56868 40236
rect 57932 39730 57988 39742
rect 57932 39678 57934 39730
rect 57986 39678 57988 39730
rect 54572 37378 54740 37380
rect 54572 37326 54574 37378
rect 54626 37326 54740 37378
rect 54572 37324 54740 37326
rect 54796 38668 55300 38724
rect 56028 39618 56084 39630
rect 56028 39566 56030 39618
rect 56082 39566 56084 39618
rect 54796 38052 54852 38668
rect 54796 37378 54852 37996
rect 55804 38050 55860 38062
rect 55804 37998 55806 38050
rect 55858 37998 55860 38050
rect 55244 37940 55300 37950
rect 55244 37938 55524 37940
rect 55244 37886 55246 37938
rect 55298 37886 55524 37938
rect 55244 37884 55524 37886
rect 55244 37874 55300 37884
rect 54796 37326 54798 37378
rect 54850 37326 54852 37378
rect 54572 37314 54628 37324
rect 54796 37314 54852 37326
rect 55468 37380 55524 37884
rect 55692 37380 55748 37390
rect 55468 37378 55748 37380
rect 55468 37326 55694 37378
rect 55746 37326 55748 37378
rect 55468 37324 55748 37326
rect 55692 37314 55748 37324
rect 54236 36654 54238 36706
rect 54290 36654 54292 36706
rect 54236 36642 54292 36654
rect 53900 36430 53902 36482
rect 53954 36430 53956 36482
rect 53900 36418 53956 36430
rect 55580 36482 55636 36494
rect 55580 36430 55582 36482
rect 55634 36430 55636 36482
rect 53788 36318 53790 36370
rect 53842 36318 53844 36370
rect 53788 36306 53844 36318
rect 54348 36372 54404 36382
rect 54404 36316 54516 36372
rect 54348 36278 54404 36316
rect 53452 35700 53508 35710
rect 53340 35698 53508 35700
rect 53340 35646 53454 35698
rect 53506 35646 53508 35698
rect 53340 35644 53508 35646
rect 53340 35252 53396 35644
rect 53452 35634 53508 35644
rect 53788 35700 53844 35710
rect 53340 35186 53396 35196
rect 52892 34860 53060 34916
rect 52780 34804 52836 34814
rect 52780 34710 52836 34748
rect 52892 34692 52948 34702
rect 52892 34598 52948 34636
rect 52556 34412 52836 34468
rect 52444 34130 52500 34188
rect 52444 34078 52446 34130
rect 52498 34078 52500 34130
rect 52444 34066 52500 34078
rect 51436 33518 51438 33570
rect 51490 33518 51492 33570
rect 51436 33506 51492 33518
rect 51884 34018 51940 34030
rect 51884 33966 51886 34018
rect 51938 33966 51940 34018
rect 50764 33460 50820 33470
rect 50764 33366 50820 33404
rect 50204 33282 50260 33292
rect 50876 33348 50932 33358
rect 49756 33236 49812 33246
rect 49644 33234 49812 33236
rect 49644 33182 49758 33234
rect 49810 33182 49812 33234
rect 49644 33180 49812 33182
rect 49644 32788 49700 33180
rect 49756 33170 49812 33180
rect 50092 33234 50148 33246
rect 50652 33236 50708 33246
rect 50092 33182 50094 33234
rect 50146 33182 50148 33234
rect 50092 33124 50148 33182
rect 50092 32788 50148 33068
rect 49644 32674 49700 32732
rect 49644 32622 49646 32674
rect 49698 32622 49700 32674
rect 49644 32610 49700 32622
rect 49756 32732 50148 32788
rect 50316 33234 50708 33236
rect 50316 33182 50654 33234
rect 50706 33182 50708 33234
rect 50316 33180 50708 33182
rect 50316 32786 50372 33180
rect 50652 33170 50708 33180
rect 50876 33234 50932 33292
rect 51884 33348 51940 33966
rect 52780 33458 52836 34412
rect 53004 34356 53060 34860
rect 53004 34242 53060 34300
rect 53788 34354 53844 35644
rect 54236 35700 54292 35710
rect 54236 35606 54292 35644
rect 54348 35586 54404 35598
rect 54348 35534 54350 35586
rect 54402 35534 54404 35586
rect 53788 34302 53790 34354
rect 53842 34302 53844 34354
rect 53788 34290 53844 34302
rect 54236 35252 54292 35262
rect 53004 34190 53006 34242
rect 53058 34190 53060 34242
rect 53004 34178 53060 34190
rect 54236 34242 54292 35196
rect 54348 34354 54404 35534
rect 54348 34302 54350 34354
rect 54402 34302 54404 34354
rect 54348 34290 54404 34302
rect 54460 34804 54516 36316
rect 55356 36260 55412 36270
rect 54684 35700 54740 35710
rect 54684 34914 54740 35644
rect 54684 34862 54686 34914
rect 54738 34862 54740 34914
rect 54684 34850 54740 34862
rect 55132 35698 55188 35710
rect 55132 35646 55134 35698
rect 55186 35646 55188 35698
rect 54460 34354 54516 34748
rect 54460 34302 54462 34354
rect 54514 34302 54516 34354
rect 54460 34290 54516 34302
rect 54236 34190 54238 34242
rect 54290 34190 54292 34242
rect 54236 34178 54292 34190
rect 55132 34244 55188 35646
rect 55356 35028 55412 36204
rect 55356 34962 55412 34972
rect 55580 34354 55636 36430
rect 55804 35476 55860 37998
rect 56028 37490 56084 39566
rect 56028 37438 56030 37490
rect 56082 37438 56084 37490
rect 56028 37426 56084 37438
rect 57708 38162 57764 38174
rect 57708 38110 57710 38162
rect 57762 38110 57764 38162
rect 56588 36260 56644 36270
rect 56588 36166 56644 36204
rect 57708 35700 57764 38110
rect 57932 37716 57988 39678
rect 57932 37650 57988 37660
rect 57708 35634 57764 35644
rect 55804 35410 55860 35420
rect 55804 34804 55860 34814
rect 55804 34710 55860 34748
rect 55580 34302 55582 34354
rect 55634 34302 55636 34354
rect 55580 34290 55636 34302
rect 55244 34244 55300 34254
rect 55132 34242 55300 34244
rect 55132 34190 55246 34242
rect 55298 34190 55300 34242
rect 55132 34188 55300 34190
rect 55244 34178 55300 34188
rect 52780 33406 52782 33458
rect 52834 33406 52836 33458
rect 52780 33394 52836 33406
rect 57932 33458 57988 33470
rect 57932 33406 57934 33458
rect 57986 33406 57988 33458
rect 51884 33282 51940 33292
rect 53004 33348 53060 33358
rect 53004 33254 53060 33292
rect 54348 33348 54404 33358
rect 50876 33182 50878 33234
rect 50930 33182 50932 33234
rect 50876 33170 50932 33182
rect 51324 33236 51380 33246
rect 51324 33142 51380 33180
rect 53676 33236 53732 33246
rect 54012 33236 54068 33246
rect 53676 33234 54068 33236
rect 53676 33182 53678 33234
rect 53730 33182 54014 33234
rect 54066 33182 54068 33234
rect 53676 33180 54068 33182
rect 53676 33170 53732 33180
rect 54012 33170 54068 33180
rect 54348 33234 54404 33292
rect 55580 33348 55636 33358
rect 55580 33254 55636 33292
rect 54348 33182 54350 33234
rect 54402 33182 54404 33234
rect 54348 33170 54404 33182
rect 51436 33124 51492 33134
rect 51436 33030 51492 33068
rect 57932 33012 57988 33406
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 57932 32946 57988 32956
rect 50556 32890 50820 32900
rect 50316 32734 50318 32786
rect 50370 32734 50372 32786
rect 49532 32498 49588 32508
rect 49756 32562 49812 32732
rect 50316 32722 50372 32734
rect 49756 32510 49758 32562
rect 49810 32510 49812 32562
rect 49196 32004 49252 32014
rect 49756 32004 49812 32510
rect 49868 32564 49924 32574
rect 49868 32470 49924 32508
rect 48972 32002 49812 32004
rect 48972 31950 49198 32002
rect 49250 31950 49812 32002
rect 48972 31948 49812 31950
rect 48860 31910 48916 31948
rect 49196 31938 49252 31948
rect 48636 31892 48692 31902
rect 48300 31890 48692 31892
rect 48300 31838 48638 31890
rect 48690 31838 48692 31890
rect 48300 31836 48692 31838
rect 48636 31826 48692 31836
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 47292 31106 47796 31108
rect 47292 31054 47294 31106
rect 47346 31054 47796 31106
rect 47292 31052 47796 31054
rect 57820 31108 57876 31118
rect 47292 31042 47348 31052
rect 57820 31014 57876 31052
rect 46732 30942 46734 30994
rect 46786 30942 46788 30994
rect 46732 30930 46788 30942
rect 58156 30994 58212 31006
rect 58156 30942 58158 30994
rect 58210 30942 58212 30994
rect 57596 30884 57652 30894
rect 58156 30884 58212 30942
rect 57596 30882 58212 30884
rect 57596 30830 57598 30882
rect 57650 30830 58212 30882
rect 57596 30828 58212 30830
rect 57596 30818 57652 30828
rect 58156 30324 58212 30828
rect 58156 30258 58212 30268
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 46396 29598 46398 29650
rect 46450 29598 46452 29650
rect 46396 29586 46452 29598
rect 43932 29362 43988 29372
rect 45612 29538 45668 29550
rect 45612 29486 45614 29538
rect 45666 29486 45668 29538
rect 43932 28084 43988 28094
rect 43932 27990 43988 28028
rect 45164 28084 45220 28094
rect 44492 27636 44548 27646
rect 44492 27542 44548 27580
rect 43036 27074 43428 27076
rect 43036 27022 43038 27074
rect 43090 27022 43428 27074
rect 43036 27020 43428 27022
rect 43484 27076 43540 27086
rect 43036 27010 43092 27020
rect 43484 26982 43540 27020
rect 45164 26514 45220 28028
rect 45612 28084 45668 29486
rect 58156 28418 58212 28430
rect 58156 28366 58158 28418
rect 58210 28366 58212 28418
rect 58156 28308 58212 28366
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 58156 28242 58212 28252
rect 50556 28186 50820 28196
rect 45612 28018 45668 28028
rect 58156 26852 58212 26862
rect 58156 26850 58324 26852
rect 58156 26798 58158 26850
rect 58210 26798 58324 26850
rect 58156 26796 58324 26798
rect 58156 26786 58212 26796
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 45164 26462 45166 26514
rect 45218 26462 45220 26514
rect 45164 26450 45220 26462
rect 58156 26402 58212 26414
rect 58156 26350 58158 26402
rect 58210 26350 58212 26402
rect 42812 26290 42868 26302
rect 42812 26238 42814 26290
rect 42866 26238 42868 26290
rect 42812 25730 42868 26238
rect 42812 25678 42814 25730
rect 42866 25678 42868 25730
rect 42812 25666 42868 25678
rect 43484 26068 43540 26078
rect 42364 25618 42756 25620
rect 42364 25566 42366 25618
rect 42418 25566 42756 25618
rect 42364 25564 42756 25566
rect 42364 25554 42420 25564
rect 42700 25508 42756 25564
rect 43372 25508 43428 25518
rect 42700 25452 42868 25508
rect 42812 25394 42868 25452
rect 42812 25342 42814 25394
rect 42866 25342 42868 25394
rect 42700 25284 42756 25294
rect 42252 24724 42308 24734
rect 42140 24722 42308 24724
rect 42140 24670 42254 24722
rect 42306 24670 42308 24722
rect 42140 24668 42308 24670
rect 41244 23938 41860 23940
rect 41244 23886 41694 23938
rect 41746 23886 41860 23938
rect 41244 23884 41860 23886
rect 42028 23938 42084 23950
rect 42028 23886 42030 23938
rect 42082 23886 42084 23938
rect 41692 23874 41748 23884
rect 40684 23716 40740 23726
rect 40684 23714 40964 23716
rect 40684 23662 40686 23714
rect 40738 23662 40964 23714
rect 40684 23660 40964 23662
rect 40684 23650 40740 23660
rect 40908 23380 40964 23660
rect 40908 23286 40964 23324
rect 40796 22148 40852 22158
rect 41132 22148 41188 23772
rect 41804 23716 41860 23726
rect 41692 23604 41748 23614
rect 40852 22092 41188 22148
rect 41244 23266 41300 23278
rect 41244 23214 41246 23266
rect 41298 23214 41300 23266
rect 41244 23044 41300 23214
rect 41692 23044 41748 23548
rect 41244 23042 41748 23044
rect 41244 22990 41694 23042
rect 41746 22990 41748 23042
rect 41244 22988 41748 22990
rect 40684 19460 40740 19470
rect 40684 19366 40740 19404
rect 40796 19012 40852 22092
rect 41132 21252 41188 21262
rect 41132 20802 41188 21196
rect 41132 20750 41134 20802
rect 41186 20750 41188 20802
rect 40908 20690 40964 20702
rect 40908 20638 40910 20690
rect 40962 20638 40964 20690
rect 40908 20356 40964 20638
rect 41132 20580 41188 20750
rect 41132 20514 41188 20524
rect 40908 20290 40964 20300
rect 41244 20188 41300 22988
rect 41692 22978 41748 22988
rect 41804 22036 41860 23660
rect 41916 23156 41972 23166
rect 42028 23156 42084 23886
rect 42140 23828 42196 24668
rect 42252 24658 42308 24668
rect 42700 24722 42756 25228
rect 42812 25172 42868 25342
rect 42924 25396 42980 25406
rect 43148 25396 43204 25406
rect 43372 25396 43428 25452
rect 42924 25394 43204 25396
rect 42924 25342 42926 25394
rect 42978 25342 43150 25394
rect 43202 25342 43204 25394
rect 42924 25340 43204 25342
rect 42924 25330 42980 25340
rect 43148 25330 43204 25340
rect 43260 25394 43428 25396
rect 43260 25342 43374 25394
rect 43426 25342 43428 25394
rect 43260 25340 43428 25342
rect 42812 25106 42868 25116
rect 43260 25060 43316 25340
rect 43372 25330 43428 25340
rect 43484 25394 43540 26012
rect 45948 26068 46004 26078
rect 45948 25974 46004 26012
rect 57932 25618 57988 25630
rect 57932 25566 57934 25618
rect 57986 25566 57988 25618
rect 43932 25508 43988 25518
rect 43932 25414 43988 25452
rect 46844 25506 46900 25518
rect 46844 25454 46846 25506
rect 46898 25454 46900 25506
rect 43484 25342 43486 25394
rect 43538 25342 43540 25394
rect 43484 25284 43540 25342
rect 43484 25218 43540 25228
rect 42700 24670 42702 24722
rect 42754 24670 42756 24722
rect 42700 24658 42756 24670
rect 43148 25004 43316 25060
rect 44828 25172 44884 25182
rect 42812 24612 42868 24622
rect 42812 24610 42980 24612
rect 42812 24558 42814 24610
rect 42866 24558 42980 24610
rect 42812 24556 42980 24558
rect 42812 24546 42868 24556
rect 42140 23762 42196 23772
rect 42252 23940 42308 23950
rect 42588 23940 42644 23950
rect 42308 23938 42644 23940
rect 42308 23886 42590 23938
rect 42642 23886 42644 23938
rect 42308 23884 42644 23886
rect 41916 23154 42084 23156
rect 41916 23102 41918 23154
rect 41970 23102 42084 23154
rect 41916 23100 42084 23102
rect 42140 23156 42196 23166
rect 42252 23156 42308 23884
rect 42588 23874 42644 23884
rect 42364 23714 42420 23726
rect 42364 23662 42366 23714
rect 42418 23662 42420 23714
rect 42364 23604 42420 23662
rect 42476 23716 42532 23726
rect 42476 23622 42532 23660
rect 42364 23538 42420 23548
rect 42700 23604 42756 23614
rect 42588 23380 42644 23390
rect 42700 23380 42756 23548
rect 42588 23378 42756 23380
rect 42588 23326 42590 23378
rect 42642 23326 42756 23378
rect 42588 23324 42756 23326
rect 42588 23314 42644 23324
rect 42140 23154 42308 23156
rect 42140 23102 42142 23154
rect 42194 23102 42308 23154
rect 42140 23100 42308 23102
rect 42812 23266 42868 23278
rect 42812 23214 42814 23266
rect 42866 23214 42868 23266
rect 41916 22260 41972 23100
rect 42140 23090 42196 23100
rect 41916 22194 41972 22204
rect 41804 21980 42308 22036
rect 41692 21812 41748 21822
rect 42140 21812 42196 21822
rect 41468 21810 42196 21812
rect 41468 21758 41694 21810
rect 41746 21758 42142 21810
rect 42194 21758 42196 21810
rect 41468 21756 42196 21758
rect 41356 20916 41412 20926
rect 41356 20802 41412 20860
rect 41356 20750 41358 20802
rect 41410 20750 41412 20802
rect 41356 20738 41412 20750
rect 41468 20692 41524 21756
rect 41692 21746 41748 21756
rect 42140 21746 42196 21756
rect 41580 21588 41636 21598
rect 41580 21494 41636 21532
rect 41692 21364 41748 21374
rect 41692 21362 41860 21364
rect 41692 21310 41694 21362
rect 41746 21310 41860 21362
rect 41692 21308 41860 21310
rect 41692 21298 41748 21308
rect 41580 20804 41636 20842
rect 41580 20738 41636 20748
rect 41692 20802 41748 20814
rect 41692 20750 41694 20802
rect 41746 20750 41748 20802
rect 41468 20626 41524 20636
rect 41580 20580 41636 20590
rect 41244 20132 41412 20188
rect 40796 18946 40852 18956
rect 41356 17668 41412 20132
rect 41580 20130 41636 20524
rect 41580 20078 41582 20130
rect 41634 20078 41636 20130
rect 41580 20066 41636 20078
rect 41692 20020 41748 20750
rect 41692 19460 41748 19964
rect 41692 19394 41748 19404
rect 41580 19012 41636 19022
rect 41636 18956 41748 19012
rect 41580 18946 41636 18956
rect 40572 17612 40852 17668
rect 40348 17500 40740 17556
rect 39116 17444 39172 17454
rect 39116 17350 39172 17388
rect 39004 16044 39172 16100
rect 38892 15986 38948 15998
rect 38892 15934 38894 15986
rect 38946 15934 38948 15986
rect 38892 15092 38948 15934
rect 39004 15874 39060 15886
rect 39004 15822 39006 15874
rect 39058 15822 39060 15874
rect 39004 15314 39060 15822
rect 39004 15262 39006 15314
rect 39058 15262 39060 15314
rect 39004 15250 39060 15262
rect 38892 15036 39060 15092
rect 38892 14530 38948 14542
rect 38892 14478 38894 14530
rect 38946 14478 38948 14530
rect 38892 13860 38948 14478
rect 39004 14532 39060 15036
rect 39004 14466 39060 14476
rect 39116 14420 39172 16044
rect 39900 16098 39956 16110
rect 39900 16046 39902 16098
rect 39954 16046 39956 16098
rect 39228 15986 39284 15998
rect 39228 15934 39230 15986
rect 39282 15934 39284 15986
rect 39228 15092 39284 15934
rect 39788 15986 39844 15998
rect 39788 15934 39790 15986
rect 39842 15934 39844 15986
rect 39788 15540 39844 15934
rect 39900 15876 39956 16046
rect 39900 15810 39956 15820
rect 40124 16100 40180 16110
rect 39788 15484 39956 15540
rect 39228 15026 39284 15036
rect 39676 15314 39732 15326
rect 39676 15262 39678 15314
rect 39730 15262 39732 15314
rect 39452 14532 39508 14542
rect 39676 14532 39732 15262
rect 39788 15314 39844 15326
rect 39788 15262 39790 15314
rect 39842 15262 39844 15314
rect 39788 15092 39844 15262
rect 39788 14642 39844 15036
rect 39788 14590 39790 14642
rect 39842 14590 39844 14642
rect 39788 14578 39844 14590
rect 39508 14476 39732 14532
rect 39452 14438 39508 14476
rect 39116 14354 39172 14364
rect 38892 13748 38948 13804
rect 39340 13860 39396 13870
rect 39340 13766 39396 13804
rect 39004 13748 39060 13758
rect 38892 13746 39060 13748
rect 38892 13694 39006 13746
rect 39058 13694 39060 13746
rect 38892 13692 39060 13694
rect 39004 13682 39060 13692
rect 38780 13580 38948 13636
rect 38444 13468 38836 13524
rect 38444 12404 38500 12414
rect 38332 12402 38500 12404
rect 38332 12350 38446 12402
rect 38498 12350 38500 12402
rect 38332 12348 38500 12350
rect 37996 11230 37998 11282
rect 38050 11230 38052 11282
rect 37996 11218 38052 11230
rect 37212 9940 37268 10556
rect 37548 11170 37604 11182
rect 38220 11172 38276 11182
rect 37548 11118 37550 11170
rect 37602 11118 37604 11170
rect 37548 10500 37604 11118
rect 38108 11170 38276 11172
rect 38108 11118 38222 11170
rect 38274 11118 38276 11170
rect 38108 11116 38276 11118
rect 38108 10836 38164 11116
rect 38220 11106 38276 11116
rect 37660 10780 38164 10836
rect 37660 10610 37716 10780
rect 37660 10558 37662 10610
rect 37714 10558 37716 10610
rect 37660 10546 37716 10558
rect 38444 10612 38500 12348
rect 38780 12402 38836 13468
rect 38780 12350 38782 12402
rect 38834 12350 38836 12402
rect 38780 11732 38836 12350
rect 38892 12180 38948 13580
rect 39900 12292 39956 15484
rect 40124 14754 40180 16044
rect 40236 15092 40292 15102
rect 40236 14998 40292 15036
rect 40124 14702 40126 14754
rect 40178 14702 40180 14754
rect 40124 14690 40180 14702
rect 39676 12236 39956 12292
rect 39116 12180 39172 12190
rect 38892 12178 39172 12180
rect 38892 12126 39118 12178
rect 39170 12126 39172 12178
rect 38892 12124 39172 12126
rect 38780 11666 38836 11676
rect 38556 10612 38612 10622
rect 38444 10610 38612 10612
rect 38444 10558 38558 10610
rect 38610 10558 38612 10610
rect 38444 10556 38612 10558
rect 37548 10434 37604 10444
rect 37884 10498 37940 10510
rect 37884 10446 37886 10498
rect 37938 10446 37940 10498
rect 37324 10388 37380 10398
rect 37884 10388 37940 10446
rect 37324 10386 37492 10388
rect 37324 10334 37326 10386
rect 37378 10334 37492 10386
rect 37324 10332 37492 10334
rect 37324 10322 37380 10332
rect 37212 9874 37268 9884
rect 37100 9202 37156 9212
rect 36988 6692 37044 6702
rect 36876 6690 37044 6692
rect 36876 6638 36990 6690
rect 37042 6638 37044 6690
rect 36876 6636 37044 6638
rect 36204 5908 36260 5918
rect 36204 5814 36260 5852
rect 36876 5908 36932 6636
rect 36988 6626 37044 6636
rect 37436 6580 37492 10332
rect 37884 10322 37940 10332
rect 38556 10276 38612 10556
rect 39004 10612 39060 10622
rect 39116 10612 39172 12124
rect 39676 12178 39732 12236
rect 39676 12126 39678 12178
rect 39730 12126 39732 12178
rect 39676 12114 39732 12126
rect 39676 11506 39732 11518
rect 39676 11454 39678 11506
rect 39730 11454 39732 11506
rect 39452 11396 39508 11406
rect 39452 11302 39508 11340
rect 39004 10610 39172 10612
rect 39004 10558 39006 10610
rect 39058 10558 39172 10610
rect 39004 10556 39172 10558
rect 39004 10546 39060 10556
rect 39452 10500 39508 10510
rect 38556 10210 38612 10220
rect 39228 10498 39508 10500
rect 39228 10446 39454 10498
rect 39506 10446 39508 10498
rect 39228 10444 39508 10446
rect 38668 9828 38724 9838
rect 38444 9714 38500 9726
rect 38444 9662 38446 9714
rect 38498 9662 38500 9714
rect 38220 9604 38276 9614
rect 38444 9604 38500 9662
rect 38556 9716 38612 9726
rect 38556 9622 38612 9660
rect 38220 9602 38500 9604
rect 38220 9550 38222 9602
rect 38274 9550 38500 9602
rect 38220 9548 38500 9550
rect 38220 8036 38276 9548
rect 38668 9042 38724 9772
rect 38780 9828 38836 9838
rect 39116 9828 39172 9838
rect 38780 9826 39172 9828
rect 38780 9774 38782 9826
rect 38834 9774 39118 9826
rect 39170 9774 39172 9826
rect 38780 9772 39172 9774
rect 38780 9762 38836 9772
rect 39116 9762 39172 9772
rect 38668 8990 38670 9042
rect 38722 8990 38724 9042
rect 38668 8978 38724 8990
rect 39116 9044 39172 9054
rect 39228 9044 39284 10444
rect 39452 10434 39508 10444
rect 39676 10500 39732 11454
rect 39788 11282 39844 12236
rect 40348 11508 40404 11518
rect 40348 11394 40404 11452
rect 40348 11342 40350 11394
rect 40402 11342 40404 11394
rect 40348 11330 40404 11342
rect 40460 11396 40516 11406
rect 40516 11340 40628 11396
rect 40460 11330 40516 11340
rect 39788 11230 39790 11282
rect 39842 11230 39844 11282
rect 39788 10724 39844 11230
rect 39788 10658 39844 10668
rect 39676 10434 39732 10444
rect 39340 10276 39396 10286
rect 39340 9826 39396 10220
rect 40460 10052 40516 10062
rect 39340 9774 39342 9826
rect 39394 9774 39396 9826
rect 39340 9762 39396 9774
rect 40012 9828 40068 9838
rect 40012 9734 40068 9772
rect 39788 9268 39844 9278
rect 39788 9174 39844 9212
rect 40460 9268 40516 9996
rect 40572 9938 40628 11340
rect 40572 9886 40574 9938
rect 40626 9886 40628 9938
rect 40572 9874 40628 9886
rect 40684 9826 40740 17500
rect 40796 16660 40852 17612
rect 40796 16594 40852 16604
rect 40908 17444 40964 17454
rect 40796 16098 40852 16110
rect 40796 16046 40798 16098
rect 40850 16046 40852 16098
rect 40796 15538 40852 16046
rect 40796 15486 40798 15538
rect 40850 15486 40852 15538
rect 40796 15474 40852 15486
rect 40908 15540 40964 17388
rect 41132 17108 41188 17118
rect 41020 16884 41076 16894
rect 41020 16790 41076 16828
rect 41020 15540 41076 15550
rect 40908 15538 41076 15540
rect 40908 15486 41022 15538
rect 41074 15486 41076 15538
rect 40908 15484 41076 15486
rect 41132 15540 41188 17052
rect 41356 16660 41412 17612
rect 41692 17666 41748 18956
rect 41692 17614 41694 17666
rect 41746 17614 41748 17666
rect 41692 17602 41748 17614
rect 41692 17332 41748 17342
rect 41580 17276 41692 17332
rect 41244 16604 41412 16660
rect 41468 16994 41524 17006
rect 41468 16942 41470 16994
rect 41522 16942 41524 16994
rect 41468 16660 41524 16942
rect 41244 16098 41300 16604
rect 41468 16594 41524 16604
rect 41356 16324 41412 16334
rect 41412 16268 41524 16324
rect 41356 16258 41412 16268
rect 41244 16046 41246 16098
rect 41298 16046 41300 16098
rect 41244 16034 41300 16046
rect 41356 16100 41412 16110
rect 41356 16006 41412 16044
rect 41468 15876 41524 16268
rect 41132 15484 41300 15540
rect 41020 15474 41076 15484
rect 41132 15314 41188 15326
rect 41132 15262 41134 15314
rect 41186 15262 41188 15314
rect 41132 14980 41188 15262
rect 41132 14914 41188 14924
rect 41132 14756 41188 14766
rect 41132 14530 41188 14700
rect 41132 14478 41134 14530
rect 41186 14478 41188 14530
rect 41132 14466 41188 14478
rect 41132 11508 41188 11518
rect 41244 11508 41300 15484
rect 41468 15204 41524 15820
rect 41580 15428 41636 17276
rect 41692 17266 41748 17276
rect 41692 17108 41748 17118
rect 41804 17108 41860 21308
rect 41916 20578 41972 20590
rect 41916 20526 41918 20578
rect 41970 20526 41972 20578
rect 41916 20244 41972 20526
rect 41916 20178 41972 20188
rect 42252 20188 42308 21980
rect 42476 21812 42532 21822
rect 42476 21718 42532 21756
rect 42812 21700 42868 23214
rect 42924 23044 42980 24556
rect 43148 24500 43204 25004
rect 43260 24836 43316 24846
rect 43260 24742 43316 24780
rect 43372 24610 43428 24622
rect 43372 24558 43374 24610
rect 43426 24558 43428 24610
rect 43148 24444 43316 24500
rect 43148 24276 43204 24286
rect 42924 22978 42980 22988
rect 43036 24164 43092 24174
rect 43036 21812 43092 24108
rect 43148 23378 43204 24220
rect 43148 23326 43150 23378
rect 43202 23326 43204 23378
rect 43148 23314 43204 23326
rect 43260 22484 43316 24444
rect 43372 24276 43428 24558
rect 43484 24500 43540 24510
rect 43484 24406 43540 24444
rect 43372 24220 43540 24276
rect 43484 24050 43540 24220
rect 43484 23998 43486 24050
rect 43538 23998 43540 24050
rect 43484 23986 43540 23998
rect 42812 21698 42980 21700
rect 42812 21646 42814 21698
rect 42866 21646 42980 21698
rect 42812 21644 42980 21646
rect 42812 21634 42868 21644
rect 42924 21252 42980 21644
rect 43036 21698 43092 21756
rect 43036 21646 43038 21698
rect 43090 21646 43092 21698
rect 43036 21634 43092 21646
rect 43148 22428 43316 22484
rect 43372 23938 43428 23950
rect 43372 23886 43374 23938
rect 43426 23886 43428 23938
rect 42924 21196 43092 21252
rect 42364 20916 42420 20926
rect 42364 20822 42420 20860
rect 42812 20804 42868 20814
rect 42588 20802 42868 20804
rect 42588 20750 42814 20802
rect 42866 20750 42868 20802
rect 42588 20748 42868 20750
rect 42588 20188 42644 20748
rect 42812 20738 42868 20748
rect 42252 20132 42644 20188
rect 42700 20580 42756 20590
rect 41916 20018 41972 20030
rect 41916 19966 41918 20018
rect 41970 19966 41972 20018
rect 41916 17892 41972 19966
rect 42252 19012 42308 20132
rect 42700 20018 42756 20524
rect 42700 19966 42702 20018
rect 42754 19966 42756 20018
rect 42700 19954 42756 19966
rect 42924 20020 42980 20030
rect 42924 19926 42980 19964
rect 42364 19012 42420 19022
rect 42252 19010 42420 19012
rect 42252 18958 42366 19010
rect 42418 18958 42420 19010
rect 42252 18956 42420 18958
rect 41916 17836 42196 17892
rect 41916 17332 41972 17836
rect 42140 17778 42196 17836
rect 42140 17726 42142 17778
rect 42194 17726 42196 17778
rect 42140 17714 42196 17726
rect 41916 17266 41972 17276
rect 41692 17106 42196 17108
rect 41692 17054 41694 17106
rect 41746 17054 42196 17106
rect 41692 17052 42196 17054
rect 41692 17042 41748 17052
rect 41804 16884 41860 16894
rect 41804 16790 41860 16828
rect 41916 16884 41972 16894
rect 41916 16882 42084 16884
rect 41916 16830 41918 16882
rect 41970 16830 42084 16882
rect 41916 16828 42084 16830
rect 41916 16772 41972 16828
rect 41916 16706 41972 16716
rect 41916 16324 41972 16334
rect 41916 16230 41972 16268
rect 42028 15986 42084 16828
rect 42028 15934 42030 15986
rect 42082 15934 42084 15986
rect 42028 15922 42084 15934
rect 41580 15372 41748 15428
rect 41580 15204 41636 15214
rect 41468 15202 41636 15204
rect 41468 15150 41582 15202
rect 41634 15150 41636 15202
rect 41468 15148 41636 15150
rect 41580 15138 41636 15148
rect 41692 14418 41748 15372
rect 42140 15314 42196 17052
rect 42140 15262 42142 15314
rect 42194 15262 42196 15314
rect 42140 15250 42196 15262
rect 42252 15986 42308 18956
rect 42364 18946 42420 18956
rect 43036 17780 43092 21196
rect 43148 20916 43204 22428
rect 43372 21700 43428 23886
rect 44268 23826 44324 23838
rect 44268 23774 44270 23826
rect 44322 23774 44324 23826
rect 44268 23268 44324 23774
rect 44268 23202 44324 23212
rect 43372 21606 43428 21644
rect 44604 23044 44660 23054
rect 43148 20188 43204 20860
rect 43260 21474 43316 21486
rect 43260 21422 43262 21474
rect 43314 21422 43316 21474
rect 43260 20802 43316 21422
rect 43708 20916 43764 20926
rect 44044 20916 44100 20926
rect 43708 20914 44044 20916
rect 43708 20862 43710 20914
rect 43762 20862 44044 20914
rect 43708 20860 44044 20862
rect 43708 20850 43764 20860
rect 44044 20822 44100 20860
rect 43260 20750 43262 20802
rect 43314 20750 43316 20802
rect 43260 20738 43316 20750
rect 44156 20578 44212 20590
rect 44156 20526 44158 20578
rect 44210 20526 44212 20578
rect 44044 20468 44100 20478
rect 43708 20244 43764 20254
rect 43932 20244 43988 20254
rect 43148 20132 43428 20188
rect 43708 20132 43876 20188
rect 42924 17724 43092 17780
rect 43260 18452 43316 18462
rect 42700 17668 42756 17678
rect 42700 17574 42756 17612
rect 42252 15934 42254 15986
rect 42306 15934 42308 15986
rect 42252 15316 42308 15934
rect 42476 16882 42532 16894
rect 42476 16830 42478 16882
rect 42530 16830 42532 16882
rect 42364 15876 42420 15886
rect 42476 15876 42532 16830
rect 42588 16884 42644 16894
rect 42588 16770 42644 16828
rect 42588 16718 42590 16770
rect 42642 16718 42644 16770
rect 42588 16706 42644 16718
rect 42420 15820 42532 15876
rect 42364 15782 42420 15820
rect 42364 15316 42420 15326
rect 42252 15260 42364 15316
rect 42364 15222 42420 15260
rect 42476 15314 42532 15820
rect 42924 15540 42980 17724
rect 43036 17556 43092 17566
rect 43260 17556 43316 18396
rect 43372 17668 43428 20132
rect 43596 19908 43652 19918
rect 43484 19234 43540 19246
rect 43484 19182 43486 19234
rect 43538 19182 43540 19234
rect 43484 18676 43540 19182
rect 43596 18900 43652 19852
rect 43708 19796 43764 19806
rect 43708 19702 43764 19740
rect 43708 19460 43764 19470
rect 43820 19460 43876 20132
rect 43708 19458 43876 19460
rect 43708 19406 43710 19458
rect 43762 19406 43876 19458
rect 43708 19404 43876 19406
rect 43708 19394 43764 19404
rect 43932 19348 43988 20188
rect 43820 19292 43988 19348
rect 44044 19346 44100 20412
rect 44156 19460 44212 20526
rect 44268 19460 44324 19470
rect 44156 19458 44324 19460
rect 44156 19406 44270 19458
rect 44322 19406 44324 19458
rect 44156 19404 44324 19406
rect 44268 19394 44324 19404
rect 44044 19294 44046 19346
rect 44098 19294 44100 19346
rect 43596 18844 43764 18900
rect 43596 18676 43652 18686
rect 43484 18674 43652 18676
rect 43484 18622 43598 18674
rect 43650 18622 43652 18674
rect 43484 18620 43652 18622
rect 43596 18610 43652 18620
rect 43596 18452 43652 18462
rect 43708 18452 43764 18844
rect 43820 18562 43876 19292
rect 44044 19282 44100 19294
rect 44044 19124 44100 19134
rect 43820 18510 43822 18562
rect 43874 18510 43876 18562
rect 43820 18498 43876 18510
rect 43932 19122 44100 19124
rect 43932 19070 44046 19122
rect 44098 19070 44100 19122
rect 43932 19068 44100 19070
rect 43596 18450 43764 18452
rect 43596 18398 43598 18450
rect 43650 18398 43764 18450
rect 43596 18396 43764 18398
rect 43596 18386 43652 18396
rect 43372 17612 43540 17668
rect 43036 17554 43260 17556
rect 43036 17502 43038 17554
rect 43090 17502 43260 17554
rect 43036 17500 43260 17502
rect 43036 17490 43092 17500
rect 43260 17462 43316 17500
rect 43372 17442 43428 17454
rect 43372 17390 43374 17442
rect 43426 17390 43428 17442
rect 43372 17108 43428 17390
rect 43372 17042 43428 17052
rect 43372 16884 43428 16894
rect 43372 16790 43428 16828
rect 42924 15484 43204 15540
rect 42476 15262 42478 15314
rect 42530 15262 42532 15314
rect 42476 15250 42532 15262
rect 43036 15316 43092 15326
rect 43036 15222 43092 15260
rect 41692 14366 41694 14418
rect 41746 14366 41748 14418
rect 41468 14306 41524 14318
rect 41468 14254 41470 14306
rect 41522 14254 41524 14306
rect 41468 14084 41524 14254
rect 41468 14018 41524 14028
rect 41692 13860 41748 14366
rect 42028 15090 42084 15102
rect 42028 15038 42030 15090
rect 42082 15038 42084 15090
rect 41804 14308 41860 14318
rect 41804 14214 41860 14252
rect 41692 13804 41860 13860
rect 41580 12738 41636 12750
rect 41580 12686 41582 12738
rect 41634 12686 41636 12738
rect 41580 12068 41636 12686
rect 41692 12068 41748 12078
rect 41580 12012 41692 12068
rect 41692 11620 41748 12012
rect 41188 11452 41300 11508
rect 41356 11564 41748 11620
rect 41804 11620 41860 13804
rect 41916 13412 41972 13422
rect 41916 12850 41972 13356
rect 42028 13188 42084 15038
rect 42140 14868 42196 14878
rect 43148 14868 43204 15484
rect 42140 14530 42196 14812
rect 43036 14812 43204 14868
rect 43484 15538 43540 17612
rect 43932 17666 43988 19068
rect 44044 19058 44100 19068
rect 44044 18564 44100 18574
rect 44044 18470 44100 18508
rect 43932 17614 43934 17666
rect 43986 17614 43988 17666
rect 43820 16996 43876 17006
rect 43820 16902 43876 16940
rect 43484 15486 43486 15538
rect 43538 15486 43540 15538
rect 43484 14868 43540 15486
rect 42140 14478 42142 14530
rect 42194 14478 42196 14530
rect 42140 13412 42196 14478
rect 42364 14756 42420 14766
rect 42364 14530 42420 14700
rect 42364 14478 42366 14530
rect 42418 14478 42420 14530
rect 42364 14466 42420 14478
rect 42252 14418 42308 14430
rect 42252 14366 42254 14418
rect 42306 14366 42308 14418
rect 42252 14084 42308 14366
rect 42812 14420 42868 14430
rect 42812 14326 42868 14364
rect 42252 14018 42308 14028
rect 43036 13412 43092 14812
rect 43484 14802 43540 14812
rect 43148 14644 43204 14654
rect 43820 14644 43876 14654
rect 43204 14588 43652 14644
rect 43148 14530 43204 14588
rect 43148 14478 43150 14530
rect 43202 14478 43204 14530
rect 43148 14466 43204 14478
rect 43260 14418 43316 14430
rect 43260 14366 43262 14418
rect 43314 14366 43316 14418
rect 43148 14308 43204 14318
rect 43260 14308 43316 14366
rect 43204 14252 43316 14308
rect 43148 14242 43204 14252
rect 43260 13746 43316 14252
rect 43484 13860 43540 13898
rect 43484 13794 43540 13804
rect 43596 13858 43652 14588
rect 43820 14550 43876 14588
rect 43932 14532 43988 17614
rect 44268 17444 44324 17454
rect 44156 14532 44212 14542
rect 43932 14530 44212 14532
rect 43932 14478 44158 14530
rect 44210 14478 44212 14530
rect 43932 14476 44212 14478
rect 43596 13806 43598 13858
rect 43650 13806 43652 13858
rect 43596 13794 43652 13806
rect 43260 13694 43262 13746
rect 43314 13694 43316 13746
rect 43260 13682 43316 13694
rect 42140 13356 42532 13412
rect 42140 13188 42196 13198
rect 42028 13186 42420 13188
rect 42028 13134 42142 13186
rect 42194 13134 42420 13186
rect 42028 13132 42420 13134
rect 42140 13122 42196 13132
rect 42028 12964 42084 12974
rect 42028 12870 42084 12908
rect 41916 12798 41918 12850
rect 41970 12798 41972 12850
rect 41916 12740 41972 12798
rect 41916 12684 42308 12740
rect 42028 11954 42084 11966
rect 42028 11902 42030 11954
rect 42082 11902 42084 11954
rect 41804 11564 41972 11620
rect 41132 11414 41188 11452
rect 41356 11284 41412 11564
rect 41804 11396 41860 11406
rect 41804 11302 41860 11340
rect 40684 9774 40686 9826
rect 40738 9774 40740 9826
rect 40684 9716 40740 9774
rect 40684 9650 40740 9660
rect 41132 11228 41412 11284
rect 40460 9174 40516 9212
rect 39116 9042 39284 9044
rect 39116 8990 39118 9042
rect 39170 8990 39284 9042
rect 39116 8988 39284 8990
rect 39340 9044 39396 9054
rect 39676 9044 39732 9054
rect 39340 9042 39732 9044
rect 39340 8990 39342 9042
rect 39394 8990 39678 9042
rect 39730 8990 39732 9042
rect 39340 8988 39732 8990
rect 38668 8148 38724 8158
rect 37324 6468 37380 6478
rect 37324 6374 37380 6412
rect 37436 6018 37492 6524
rect 37436 5966 37438 6018
rect 37490 5966 37492 6018
rect 37436 5954 37492 5966
rect 37996 7980 38276 8036
rect 38556 8146 38724 8148
rect 38556 8094 38670 8146
rect 38722 8094 38724 8146
rect 38556 8092 38724 8094
rect 36876 5842 36932 5852
rect 37660 5796 37716 5806
rect 37660 5702 37716 5740
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35644 5012 35700 5022
rect 35644 4918 35700 4956
rect 35084 4898 35140 4910
rect 35084 4846 35086 4898
rect 35138 4846 35140 4898
rect 35084 4564 35140 4846
rect 35084 4498 35140 4508
rect 35308 4898 35364 4910
rect 35308 4846 35310 4898
rect 35362 4846 35364 4898
rect 35308 4452 35364 4846
rect 35532 4898 35588 4910
rect 35532 4846 35534 4898
rect 35586 4846 35588 4898
rect 35532 4564 35588 4846
rect 37884 4788 37940 4798
rect 37996 4788 38052 7980
rect 38556 6802 38612 8092
rect 38668 8082 38724 8092
rect 38780 8036 38836 8046
rect 38780 8034 38948 8036
rect 38780 7982 38782 8034
rect 38834 7982 38948 8034
rect 38780 7980 38948 7982
rect 38780 7970 38836 7980
rect 38892 7252 38948 7980
rect 39004 8034 39060 8046
rect 39004 7982 39006 8034
rect 39058 7982 39060 8034
rect 39004 7476 39060 7982
rect 39116 8036 39172 8988
rect 39340 8978 39396 8988
rect 39676 8978 39732 8988
rect 39788 8818 39844 8830
rect 39788 8766 39790 8818
rect 39842 8766 39844 8818
rect 39788 8428 39844 8766
rect 39788 8372 39956 8428
rect 39116 7970 39172 7980
rect 39004 7410 39060 7420
rect 38892 7196 39172 7252
rect 39116 6914 39172 7196
rect 39116 6862 39118 6914
rect 39170 6862 39172 6914
rect 39116 6850 39172 6862
rect 38556 6750 38558 6802
rect 38610 6750 38612 6802
rect 38556 6738 38612 6750
rect 38108 6692 38164 6702
rect 38668 6692 38724 6702
rect 39004 6692 39060 6702
rect 38164 6636 38388 6692
rect 38108 6598 38164 6636
rect 38332 5908 38388 6636
rect 38724 6690 39060 6692
rect 38724 6638 39006 6690
rect 39058 6638 39060 6690
rect 38724 6636 39060 6638
rect 38668 6598 38724 6636
rect 39004 6626 39060 6636
rect 38444 6468 38500 6478
rect 39116 6468 39172 6478
rect 38500 6466 39172 6468
rect 38500 6414 39118 6466
rect 39170 6414 39172 6466
rect 38500 6412 39172 6414
rect 38444 6374 38500 6412
rect 38444 5908 38500 5918
rect 38332 5852 38444 5908
rect 38444 5814 38500 5852
rect 38332 5682 38388 5694
rect 38332 5630 38334 5682
rect 38386 5630 38388 5682
rect 38332 5124 38388 5630
rect 38444 5124 38500 5134
rect 38332 5122 38500 5124
rect 38332 5070 38446 5122
rect 38498 5070 38500 5122
rect 38332 5068 38500 5070
rect 37940 4732 38052 4788
rect 37884 4722 37940 4732
rect 35532 4498 35588 4508
rect 38444 4564 38500 5068
rect 38668 5124 38724 5134
rect 38668 5030 38724 5068
rect 39004 5124 39060 6412
rect 39116 6402 39172 6412
rect 39900 6132 39956 8372
rect 39116 6130 39956 6132
rect 39116 6078 39902 6130
rect 39954 6078 39956 6130
rect 39116 6076 39956 6078
rect 39116 5906 39172 6076
rect 39900 6066 39956 6076
rect 39116 5854 39118 5906
rect 39170 5854 39172 5906
rect 39116 5842 39172 5854
rect 39676 5908 39732 5918
rect 39676 5814 39732 5852
rect 40012 5908 40068 5918
rect 39452 5796 39508 5806
rect 40012 5796 40068 5852
rect 39452 5348 39508 5740
rect 39900 5794 40068 5796
rect 39900 5742 40014 5794
rect 40066 5742 40068 5794
rect 39900 5740 40068 5742
rect 39788 5572 39844 5582
rect 39004 5058 39060 5068
rect 39116 5236 39172 5246
rect 38892 5012 38948 5022
rect 38444 4498 38500 4508
rect 38780 5010 38948 5012
rect 38780 4958 38894 5010
rect 38946 4958 38948 5010
rect 38780 4956 38948 4958
rect 35084 4340 35140 4350
rect 35028 4338 35140 4340
rect 35028 4286 35086 4338
rect 35138 4286 35140 4338
rect 35028 4284 35140 4286
rect 34972 4246 35028 4284
rect 35084 4274 35140 4284
rect 34412 4228 34468 4238
rect 34412 4134 34468 4172
rect 35308 4226 35364 4396
rect 38556 4340 38612 4350
rect 38780 4340 38836 4956
rect 38892 4946 38948 4956
rect 39004 4452 39060 4462
rect 39004 4358 39060 4396
rect 38556 4338 38836 4340
rect 38556 4286 38558 4338
rect 38610 4286 38836 4338
rect 38556 4284 38836 4286
rect 38556 4274 38612 4284
rect 35308 4174 35310 4226
rect 35362 4174 35364 4226
rect 35308 4162 35364 4174
rect 38108 4228 38164 4238
rect 38164 4172 38500 4228
rect 38108 4134 38164 4172
rect 32956 3614 32958 3666
rect 33010 3614 33012 3666
rect 32956 3602 33012 3614
rect 33068 4060 33572 4116
rect 35868 4116 35924 4126
rect 32172 3556 32228 3566
rect 31836 3554 32228 3556
rect 31836 3502 32174 3554
rect 32226 3502 32228 3554
rect 31836 3500 32228 3502
rect 32172 3490 32228 3500
rect 33068 3554 33124 4060
rect 35868 4022 35924 4060
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 33068 3502 33070 3554
rect 33122 3502 33124 3554
rect 33068 3490 33124 3502
rect 38444 3556 38500 4172
rect 38556 3556 38612 3566
rect 38444 3554 38612 3556
rect 38444 3502 38558 3554
rect 38610 3502 38612 3554
rect 38444 3500 38612 3502
rect 38556 3490 38612 3500
rect 38668 3442 38724 4284
rect 38892 3556 38948 3566
rect 39116 3556 39172 5180
rect 39340 5124 39396 5134
rect 39340 4450 39396 5068
rect 39452 5122 39508 5292
rect 39452 5070 39454 5122
rect 39506 5070 39508 5122
rect 39452 5058 39508 5070
rect 39676 5348 39732 5358
rect 39788 5348 39844 5516
rect 39676 5346 39844 5348
rect 39676 5294 39678 5346
rect 39730 5294 39844 5346
rect 39676 5292 39844 5294
rect 39900 5346 39956 5740
rect 40012 5730 40068 5740
rect 40348 5908 40404 5918
rect 39900 5294 39902 5346
rect 39954 5294 39956 5346
rect 39564 4564 39620 4574
rect 39564 4470 39620 4508
rect 39340 4398 39342 4450
rect 39394 4398 39396 4450
rect 39340 4386 39396 4398
rect 39676 4226 39732 5292
rect 39900 5282 39956 5294
rect 40012 5460 40068 5470
rect 40012 5010 40068 5404
rect 40348 5234 40404 5852
rect 40796 5906 40852 5918
rect 40796 5854 40798 5906
rect 40850 5854 40852 5906
rect 40572 5572 40628 5582
rect 40572 5346 40628 5516
rect 40572 5294 40574 5346
rect 40626 5294 40628 5346
rect 40572 5282 40628 5294
rect 40796 5348 40852 5854
rect 40796 5254 40852 5292
rect 40348 5182 40350 5234
rect 40402 5182 40404 5234
rect 40348 5170 40404 5182
rect 40012 4958 40014 5010
rect 40066 4958 40068 5010
rect 40012 4946 40068 4958
rect 40460 5124 40516 5134
rect 40460 4676 40516 5068
rect 40460 4610 40516 4620
rect 39676 4174 39678 4226
rect 39730 4174 39732 4226
rect 39676 4162 39732 4174
rect 38892 3554 39172 3556
rect 38892 3502 38894 3554
rect 38946 3502 39172 3554
rect 38892 3500 39172 3502
rect 38892 3490 38948 3500
rect 38668 3390 38670 3442
rect 38722 3390 38724 3442
rect 38668 3378 38724 3390
rect 41132 3332 41188 11228
rect 41468 11170 41524 11182
rect 41468 11118 41470 11170
rect 41522 11118 41524 11170
rect 41468 10836 41524 11118
rect 41468 10770 41524 10780
rect 41692 11172 41748 11182
rect 41244 10498 41300 10510
rect 41244 10446 41246 10498
rect 41298 10446 41300 10498
rect 41244 10386 41300 10446
rect 41244 10334 41246 10386
rect 41298 10334 41300 10386
rect 41244 7364 41300 10334
rect 41692 10498 41748 11116
rect 41692 10446 41694 10498
rect 41746 10446 41748 10498
rect 41692 10386 41748 10446
rect 41692 10334 41694 10386
rect 41746 10334 41748 10386
rect 41692 10322 41748 10334
rect 41356 9716 41412 9726
rect 41356 9622 41412 9660
rect 41804 9044 41860 9054
rect 41916 9044 41972 11564
rect 42028 11396 42084 11902
rect 42028 11330 42084 11340
rect 42252 11394 42308 12684
rect 42364 12178 42420 13132
rect 42364 12126 42366 12178
rect 42418 12126 42420 12178
rect 42364 12114 42420 12126
rect 42252 11342 42254 11394
rect 42306 11342 42308 11394
rect 42252 11284 42308 11342
rect 42252 11218 42308 11228
rect 42364 11170 42420 11182
rect 42364 11118 42366 11170
rect 42418 11118 42420 11170
rect 42140 10948 42196 10958
rect 42140 10610 42196 10892
rect 42140 10558 42142 10610
rect 42194 10558 42196 10610
rect 42140 10546 42196 10558
rect 42364 10612 42420 11118
rect 42364 10518 42420 10556
rect 42476 10388 42532 13356
rect 43036 13346 43092 13356
rect 43484 13636 43540 13646
rect 43484 13074 43540 13580
rect 43484 13022 43486 13074
rect 43538 13022 43540 13074
rect 43484 13010 43540 13022
rect 42588 12964 42644 12974
rect 42588 12870 42644 12908
rect 42812 12962 42868 12974
rect 42812 12910 42814 12962
rect 42866 12910 42868 12962
rect 42588 12068 42644 12078
rect 42812 12068 42868 12910
rect 42644 12012 42868 12068
rect 42924 12180 42980 12190
rect 42588 11974 42644 12012
rect 42924 11282 42980 12124
rect 43372 12180 43428 12190
rect 43372 12086 43428 12124
rect 43596 12066 43652 12078
rect 43596 12014 43598 12066
rect 43650 12014 43652 12066
rect 43596 11788 43652 12014
rect 44044 12068 44100 12078
rect 44044 11974 44100 12012
rect 43596 11732 43876 11788
rect 43820 11506 43876 11732
rect 43820 11454 43822 11506
rect 43874 11454 43876 11506
rect 43820 11442 43876 11454
rect 43372 11396 43428 11406
rect 43372 11302 43428 11340
rect 43708 11396 43764 11406
rect 43708 11302 43764 11340
rect 42924 11230 42926 11282
rect 42978 11230 42980 11282
rect 42924 11172 42980 11230
rect 43932 11284 43988 11294
rect 43932 11190 43988 11228
rect 42924 11106 42980 11116
rect 44156 11060 44212 14476
rect 43932 11004 44212 11060
rect 43036 10612 43092 10622
rect 43036 10518 43092 10556
rect 41804 9042 41972 9044
rect 41804 8990 41806 9042
rect 41858 8990 41972 9042
rect 41804 8988 41972 8990
rect 41804 8978 41860 8988
rect 41244 7298 41300 7308
rect 41468 8260 41524 8270
rect 41468 6356 41524 8204
rect 41916 8258 41972 8988
rect 42252 10332 42532 10388
rect 42252 9042 42308 10332
rect 43820 9828 43876 9838
rect 42252 8990 42254 9042
rect 42306 8990 42308 9042
rect 42252 8428 42308 8990
rect 41916 8206 41918 8258
rect 41970 8206 41972 8258
rect 41916 8194 41972 8206
rect 42028 8372 42308 8428
rect 42588 9716 42644 9726
rect 42588 9154 42644 9660
rect 43820 9602 43876 9772
rect 43820 9550 43822 9602
rect 43874 9550 43876 9602
rect 42588 9102 42590 9154
rect 42642 9102 42644 9154
rect 42028 7700 42084 8372
rect 42476 8260 42532 8270
rect 42476 8166 42532 8204
rect 42588 8258 42644 9102
rect 42924 9100 43204 9156
rect 42812 9042 42868 9054
rect 42812 8990 42814 9042
rect 42866 8990 42868 9042
rect 42812 8372 42868 8990
rect 42812 8306 42868 8316
rect 42588 8206 42590 8258
rect 42642 8206 42644 8258
rect 42588 8194 42644 8206
rect 42700 8148 42756 8158
rect 42924 8148 42980 9100
rect 43148 9042 43204 9100
rect 43148 8990 43150 9042
rect 43202 8990 43204 9042
rect 43148 8978 43204 8990
rect 43820 9044 43876 9550
rect 43820 8978 43876 8988
rect 43036 8930 43092 8942
rect 43036 8878 43038 8930
rect 43090 8878 43092 8930
rect 43036 8260 43092 8878
rect 43148 8372 43204 8382
rect 43148 8278 43204 8316
rect 43932 8372 43988 11004
rect 44268 10948 44324 17388
rect 44604 16996 44660 22988
rect 44716 20018 44772 20030
rect 44716 19966 44718 20018
rect 44770 19966 44772 20018
rect 44716 18564 44772 19966
rect 44716 18498 44772 18508
rect 44604 16930 44660 16940
rect 44828 15540 44884 25116
rect 46844 24834 46900 25454
rect 47068 25508 47124 25518
rect 47068 25394 47124 25452
rect 55580 25508 55636 25518
rect 55580 25414 55636 25452
rect 47068 25342 47070 25394
rect 47122 25342 47124 25394
rect 47068 25330 47124 25342
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 57932 24948 57988 25566
rect 58156 25620 58212 26350
rect 58268 26292 58324 26796
rect 58268 26226 58324 26236
rect 58156 25554 58212 25564
rect 57932 24882 57988 24892
rect 46844 24782 46846 24834
rect 46898 24782 46900 24834
rect 46844 24770 46900 24782
rect 46172 24722 46228 24734
rect 46172 24670 46174 24722
rect 46226 24670 46228 24722
rect 46172 24500 46228 24670
rect 46620 24722 46676 24734
rect 46620 24670 46622 24722
rect 46674 24670 46676 24722
rect 46228 24444 46452 24500
rect 46172 24434 46228 24444
rect 45836 24052 45892 24062
rect 45836 24050 46116 24052
rect 45836 23998 45838 24050
rect 45890 23998 46116 24050
rect 45836 23996 46116 23998
rect 45836 23986 45892 23996
rect 45948 23826 46004 23838
rect 45948 23774 45950 23826
rect 46002 23774 46004 23826
rect 45500 23716 45556 23726
rect 45500 23622 45556 23660
rect 45724 23714 45780 23726
rect 45724 23662 45726 23714
rect 45778 23662 45780 23714
rect 44940 23268 44996 23278
rect 44940 23174 44996 23212
rect 45388 23154 45444 23166
rect 45388 23102 45390 23154
rect 45442 23102 45444 23154
rect 45388 23044 45444 23102
rect 45388 22978 45444 22988
rect 45052 22930 45108 22942
rect 45052 22878 45054 22930
rect 45106 22878 45108 22930
rect 44940 22372 44996 22382
rect 44940 22278 44996 22316
rect 45052 22260 45108 22878
rect 45500 22932 45556 22942
rect 45724 22932 45780 23662
rect 45948 23604 46004 23774
rect 46060 23828 46116 23996
rect 46396 24050 46452 24444
rect 46620 24164 46676 24670
rect 46396 23998 46398 24050
rect 46450 23998 46452 24050
rect 46396 23986 46452 23998
rect 46508 24162 46676 24164
rect 46508 24110 46622 24162
rect 46674 24110 46676 24162
rect 46508 24108 46676 24110
rect 46508 23828 46564 24108
rect 46620 24098 46676 24108
rect 46956 24164 47012 24174
rect 47516 24164 47572 24174
rect 46956 24162 47572 24164
rect 46956 24110 46958 24162
rect 47010 24110 47518 24162
rect 47570 24110 47572 24162
rect 46956 24108 47572 24110
rect 46956 24098 47012 24108
rect 47516 24098 47572 24108
rect 57932 24050 57988 24062
rect 57932 23998 57934 24050
rect 57986 23998 57988 24050
rect 46060 23772 46564 23828
rect 47292 23938 47348 23950
rect 47292 23886 47294 23938
rect 47346 23886 47348 23938
rect 45948 23538 46004 23548
rect 47292 23604 47348 23886
rect 50092 23940 50148 23950
rect 50092 23826 50148 23884
rect 55580 23940 55636 23950
rect 55580 23846 55636 23884
rect 50092 23774 50094 23826
rect 50146 23774 50148 23826
rect 50092 23762 50148 23774
rect 47292 23538 47348 23548
rect 47852 23714 47908 23726
rect 47852 23662 47854 23714
rect 47906 23662 47908 23714
rect 46172 23268 46228 23278
rect 46172 23154 46228 23212
rect 46172 23102 46174 23154
rect 46226 23102 46228 23154
rect 46172 23090 46228 23102
rect 47852 23156 47908 23662
rect 49756 23714 49812 23726
rect 49756 23662 49758 23714
rect 49810 23662 49812 23714
rect 49756 23266 49812 23662
rect 57932 23604 57988 23998
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 57932 23538 57988 23548
rect 50556 23482 50820 23492
rect 49756 23214 49758 23266
rect 49810 23214 49812 23266
rect 49756 23202 49812 23214
rect 47852 23090 47908 23100
rect 48748 23156 48804 23166
rect 45500 22930 45780 22932
rect 45500 22878 45502 22930
rect 45554 22878 45780 22930
rect 45500 22876 45780 22878
rect 46396 23042 46452 23054
rect 46396 22990 46398 23042
rect 46450 22990 46452 23042
rect 45276 22484 45332 22494
rect 45276 22370 45332 22428
rect 45276 22318 45278 22370
rect 45330 22318 45332 22370
rect 45276 22306 45332 22318
rect 45052 22194 45108 22204
rect 45500 22146 45556 22876
rect 45612 22596 45668 22606
rect 46396 22596 46452 22990
rect 46844 23044 46900 23054
rect 46844 22950 46900 22988
rect 45612 22594 46452 22596
rect 45612 22542 45614 22594
rect 45666 22542 46452 22594
rect 45612 22540 46452 22542
rect 45612 22530 45668 22540
rect 45724 22372 45780 22382
rect 45724 22278 45780 22316
rect 46396 22370 46452 22540
rect 48748 22484 48804 23100
rect 49084 23156 49140 23166
rect 49084 23062 49140 23100
rect 48860 23044 48916 23054
rect 48916 22988 49028 23044
rect 48860 22950 48916 22988
rect 48972 22820 49028 22988
rect 48972 22764 49252 22820
rect 49196 22594 49252 22764
rect 49196 22542 49198 22594
rect 49250 22542 49252 22594
rect 49196 22530 49252 22542
rect 48972 22484 49028 22494
rect 48748 22482 49028 22484
rect 48748 22430 48974 22482
rect 49026 22430 49028 22482
rect 48748 22428 49028 22430
rect 48972 22418 49028 22428
rect 57932 22482 57988 22494
rect 57932 22430 57934 22482
rect 57986 22430 57988 22482
rect 46396 22318 46398 22370
rect 46450 22318 46452 22370
rect 46396 22306 46452 22318
rect 51100 22372 51156 22382
rect 46172 22260 46228 22270
rect 46172 22166 46228 22204
rect 45500 22094 45502 22146
rect 45554 22094 45556 22146
rect 44940 20244 44996 20254
rect 44940 20018 44996 20188
rect 44940 19966 44942 20018
rect 44994 19966 44996 20018
rect 44940 19954 44996 19966
rect 45500 18452 45556 22094
rect 46284 22146 46340 22158
rect 46284 22094 46286 22146
rect 46338 22094 46340 22146
rect 46284 21140 46340 22094
rect 49532 22148 49588 22158
rect 49532 22146 49812 22148
rect 49532 22094 49534 22146
rect 49586 22094 49812 22146
rect 49532 22092 49812 22094
rect 49532 22082 49588 22092
rect 49756 21586 49812 22092
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 51100 21810 51156 22316
rect 55580 22372 55636 22382
rect 55580 22278 55636 22316
rect 51100 21758 51102 21810
rect 51154 21758 51156 21810
rect 51100 21746 51156 21758
rect 49756 21534 49758 21586
rect 49810 21534 49812 21586
rect 49532 21474 49588 21486
rect 49532 21422 49534 21474
rect 49586 21422 49588 21474
rect 46060 21084 46788 21140
rect 45612 20690 45668 20702
rect 45612 20638 45614 20690
rect 45666 20638 45668 20690
rect 45612 20468 45668 20638
rect 46060 20690 46116 21084
rect 46060 20638 46062 20690
rect 46114 20638 46116 20690
rect 46060 20626 46116 20638
rect 46172 20692 46228 20702
rect 46172 20598 46228 20636
rect 46732 20690 46788 21084
rect 47292 20916 47348 20926
rect 46732 20638 46734 20690
rect 46786 20638 46788 20690
rect 46732 20626 46788 20638
rect 46956 20804 47012 20814
rect 45612 20402 45668 20412
rect 45836 20578 45892 20590
rect 45836 20526 45838 20578
rect 45890 20526 45892 20578
rect 45836 20188 45892 20526
rect 45836 20132 46004 20188
rect 45948 20066 46004 20076
rect 46172 20132 46228 20142
rect 46732 20132 46788 20142
rect 46172 20130 46788 20132
rect 46172 20078 46174 20130
rect 46226 20078 46734 20130
rect 46786 20078 46788 20130
rect 46172 20076 46788 20078
rect 46172 20066 46228 20076
rect 46060 20018 46116 20030
rect 46060 19966 46062 20018
rect 46114 19966 46116 20018
rect 45948 19908 46004 19918
rect 45948 19814 46004 19852
rect 45836 18452 45892 18462
rect 45500 18450 45892 18452
rect 45500 18398 45838 18450
rect 45890 18398 45892 18450
rect 45500 18396 45892 18398
rect 45724 17666 45780 17678
rect 45724 17614 45726 17666
rect 45778 17614 45780 17666
rect 45724 16882 45780 17614
rect 45724 16830 45726 16882
rect 45778 16830 45780 16882
rect 45388 16324 45444 16334
rect 45052 15540 45108 15550
rect 44828 15538 45332 15540
rect 44828 15486 45054 15538
rect 45106 15486 45332 15538
rect 44828 15484 45332 15486
rect 45052 15474 45108 15484
rect 45276 14532 45332 15484
rect 45388 15426 45444 16268
rect 45724 16212 45780 16830
rect 45724 16146 45780 16156
rect 45836 15538 45892 18396
rect 46060 18452 46116 19966
rect 46284 19796 46340 19806
rect 46284 19234 46340 19740
rect 46284 19182 46286 19234
rect 46338 19182 46340 19234
rect 46284 19170 46340 19182
rect 46620 19236 46676 19246
rect 46732 19236 46788 20076
rect 46620 19234 46788 19236
rect 46620 19182 46622 19234
rect 46674 19182 46788 19234
rect 46620 19180 46788 19182
rect 46844 20018 46900 20030
rect 46844 19966 46846 20018
rect 46898 19966 46900 20018
rect 46620 19170 46676 19180
rect 46844 19012 46900 19966
rect 46956 19458 47012 20748
rect 47292 20802 47348 20860
rect 48636 20916 48692 20926
rect 48636 20822 48692 20860
rect 49532 20916 49588 21422
rect 49532 20822 49588 20860
rect 47292 20750 47294 20802
rect 47346 20750 47348 20802
rect 47292 20188 47348 20750
rect 47964 20804 48020 20814
rect 47964 20710 48020 20748
rect 48860 20802 48916 20814
rect 48860 20750 48862 20802
rect 48914 20750 48916 20802
rect 48860 20692 48916 20750
rect 49756 20802 49812 21534
rect 50428 21588 50484 21598
rect 50764 21588 50820 21598
rect 50428 21586 50820 21588
rect 50428 21534 50430 21586
rect 50482 21534 50766 21586
rect 50818 21534 50820 21586
rect 50428 21532 50820 21534
rect 50428 21522 50484 21532
rect 50764 21522 50820 21532
rect 57932 21588 57988 22430
rect 58156 22260 58212 22270
rect 58156 21810 58212 22204
rect 58156 21758 58158 21810
rect 58210 21758 58212 21810
rect 58156 21746 58212 21758
rect 57932 21522 57988 21532
rect 49756 20750 49758 20802
rect 49810 20750 49812 20802
rect 49756 20738 49812 20750
rect 48860 20626 48916 20636
rect 50316 20690 50372 20702
rect 50316 20638 50318 20690
rect 50370 20638 50372 20690
rect 50316 20188 50372 20638
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 58156 20244 58212 20282
rect 47068 20132 47124 20142
rect 47292 20132 47572 20188
rect 47068 19794 47124 20076
rect 47516 20018 47572 20132
rect 49196 20132 49252 20142
rect 47516 19966 47518 20018
rect 47570 19966 47572 20018
rect 47516 19954 47572 19966
rect 47964 20018 48020 20030
rect 47964 19966 47966 20018
rect 48018 19966 48020 20018
rect 47068 19742 47070 19794
rect 47122 19742 47124 19794
rect 47068 19730 47124 19742
rect 47964 19796 48020 19966
rect 47964 19730 48020 19740
rect 48972 19796 49028 19806
rect 46956 19406 46958 19458
rect 47010 19406 47012 19458
rect 46956 19394 47012 19406
rect 48972 19346 49028 19740
rect 49196 19458 49252 20076
rect 49308 20130 49364 20142
rect 50316 20132 50484 20188
rect 58156 20178 58212 20188
rect 49308 20078 49310 20130
rect 49362 20078 49364 20130
rect 49308 19796 49364 20078
rect 49308 19730 49364 19740
rect 49532 20018 49588 20030
rect 49532 19966 49534 20018
rect 49586 19966 49588 20018
rect 49532 19684 49588 19966
rect 49532 19628 49812 19684
rect 49196 19406 49198 19458
rect 49250 19406 49252 19458
rect 49196 19394 49252 19406
rect 48972 19294 48974 19346
rect 49026 19294 49028 19346
rect 48972 19282 49028 19294
rect 49532 19124 49588 19134
rect 49532 19030 49588 19068
rect 46060 18386 46116 18396
rect 46732 19010 46900 19012
rect 46732 18958 46846 19010
rect 46898 18958 46900 19010
rect 46732 18956 46900 18958
rect 45948 18340 46004 18350
rect 45948 17778 46004 18284
rect 45948 17726 45950 17778
rect 46002 17726 46004 17778
rect 45948 16770 46004 17726
rect 45948 16718 45950 16770
rect 46002 16718 46004 16770
rect 45948 16706 46004 16718
rect 46284 18340 46340 18350
rect 46732 18340 46788 18956
rect 46844 18946 46900 18956
rect 49756 18562 49812 19628
rect 49756 18510 49758 18562
rect 49810 18510 49812 18562
rect 49756 18498 49812 18510
rect 50092 19346 50148 19358
rect 50092 19294 50094 19346
rect 50146 19294 50148 19346
rect 48748 18452 48804 18462
rect 46284 18338 46788 18340
rect 46284 18286 46286 18338
rect 46338 18286 46788 18338
rect 46284 18284 46788 18286
rect 46844 18338 46900 18350
rect 46844 18286 46846 18338
rect 46898 18286 46900 18338
rect 45836 15486 45838 15538
rect 45890 15486 45892 15538
rect 45836 15474 45892 15486
rect 45388 15374 45390 15426
rect 45442 15374 45444 15426
rect 45388 15362 45444 15374
rect 45612 15314 45668 15326
rect 45612 15262 45614 15314
rect 45666 15262 45668 15314
rect 45612 15092 45668 15262
rect 45948 15316 46004 15326
rect 45388 14532 45444 14542
rect 45276 14530 45444 14532
rect 45276 14478 45390 14530
rect 45442 14478 45444 14530
rect 45276 14476 45444 14478
rect 45052 14420 45108 14430
rect 44828 14306 44884 14318
rect 44828 14254 44830 14306
rect 44882 14254 44884 14306
rect 44828 13860 44884 14254
rect 44940 14308 44996 14318
rect 44940 14214 44996 14252
rect 44940 13972 44996 13982
rect 45052 13972 45108 14364
rect 44940 13970 45108 13972
rect 44940 13918 44942 13970
rect 44994 13918 45108 13970
rect 44940 13916 45108 13918
rect 45164 13972 45220 13982
rect 44940 13906 44996 13916
rect 45164 13878 45220 13916
rect 44828 13766 44884 13804
rect 45276 13412 45332 14476
rect 45388 14466 45444 14476
rect 45500 13860 45556 13870
rect 45500 13766 45556 13804
rect 45388 13636 45444 13646
rect 45388 13542 45444 13580
rect 45612 13524 45668 15036
rect 45836 15202 45892 15214
rect 45836 15150 45838 15202
rect 45890 15150 45892 15202
rect 45836 14868 45892 15150
rect 45836 14802 45892 14812
rect 45836 14644 45892 14654
rect 45948 14644 46004 15260
rect 45836 14642 46004 14644
rect 45836 14590 45838 14642
rect 45890 14590 46004 14642
rect 45836 14588 46004 14590
rect 46172 15314 46228 15326
rect 46172 15262 46174 15314
rect 46226 15262 46228 15314
rect 46172 14644 46228 15262
rect 45836 14578 45892 14588
rect 46172 14578 46228 14588
rect 45724 14308 45780 14318
rect 45724 14214 45780 14252
rect 45948 14306 46004 14318
rect 45948 14254 45950 14306
rect 46002 14254 46004 14306
rect 45836 13748 45892 13758
rect 45948 13748 46004 14254
rect 45892 13692 46004 13748
rect 46172 14308 46228 14318
rect 45836 13654 45892 13692
rect 46172 13636 46228 14252
rect 46172 13570 46228 13580
rect 45612 13458 45668 13468
rect 46284 13412 46340 18284
rect 46508 17668 46564 17678
rect 46508 17574 46564 17612
rect 46844 17554 46900 18286
rect 47516 18338 47572 18350
rect 47516 18286 47518 18338
rect 47570 18286 47572 18338
rect 47404 18228 47460 18238
rect 47292 18226 47460 18228
rect 47292 18174 47406 18226
rect 47458 18174 47460 18226
rect 47292 18172 47460 18174
rect 47068 17668 47124 17678
rect 47068 17574 47124 17612
rect 47292 17668 47348 18172
rect 47404 18162 47460 18172
rect 46844 17502 46846 17554
rect 46898 17502 46900 17554
rect 46844 16996 46900 17502
rect 46844 16930 46900 16940
rect 46956 17556 47012 17566
rect 46956 16882 47012 17500
rect 46956 16830 46958 16882
rect 47010 16830 47012 16882
rect 46956 16818 47012 16830
rect 47180 16884 47236 16894
rect 47292 16884 47348 17612
rect 47516 17780 47572 18286
rect 47404 17556 47460 17566
rect 47404 17442 47460 17500
rect 47404 17390 47406 17442
rect 47458 17390 47460 17442
rect 47404 17378 47460 17390
rect 47180 16882 47348 16884
rect 47180 16830 47182 16882
rect 47234 16830 47348 16882
rect 47180 16828 47348 16830
rect 47516 16884 47572 17724
rect 48748 17778 48804 18396
rect 49644 18452 49700 18462
rect 49644 18358 49700 18396
rect 48748 17726 48750 17778
rect 48802 17726 48804 17778
rect 48748 17714 48804 17726
rect 49532 17780 49588 17790
rect 48076 17668 48132 17678
rect 48076 17574 48132 17612
rect 48636 17668 48692 17678
rect 48636 17574 48692 17612
rect 49196 17668 49252 17678
rect 49196 17574 49252 17612
rect 49532 17666 49588 17724
rect 49532 17614 49534 17666
rect 49586 17614 49588 17666
rect 49532 17602 49588 17614
rect 50092 17556 50148 19294
rect 50428 19236 50484 20132
rect 50092 17490 50148 17500
rect 50204 19124 50260 19134
rect 50204 17668 50260 19068
rect 50428 18452 50484 19180
rect 51436 19236 51492 19246
rect 51436 19142 51492 19180
rect 52108 19124 52164 19134
rect 52668 19124 52724 19134
rect 52108 19122 52724 19124
rect 52108 19070 52110 19122
rect 52162 19070 52670 19122
rect 52722 19070 52724 19122
rect 52108 19068 52724 19070
rect 52108 19058 52164 19068
rect 52668 19058 52724 19068
rect 53004 19010 53060 19022
rect 53004 18958 53006 19010
rect 53058 18958 53060 19010
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 50540 18452 50596 18462
rect 50428 18450 50596 18452
rect 50428 18398 50542 18450
rect 50594 18398 50596 18450
rect 50428 18396 50596 18398
rect 50540 18386 50596 18396
rect 50316 18340 50372 18350
rect 50316 18246 50372 18284
rect 51660 18340 51716 18350
rect 50204 16994 50260 17612
rect 51324 17668 51380 17678
rect 51324 17574 51380 17612
rect 50652 17556 50708 17566
rect 50652 17462 50708 17500
rect 51100 17556 51156 17566
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 50204 16942 50206 16994
rect 50258 16942 50260 16994
rect 50204 16930 50260 16942
rect 47180 16818 47236 16828
rect 47516 16818 47572 16828
rect 51100 16882 51156 17500
rect 51660 17554 51716 18284
rect 53004 17668 53060 18958
rect 58156 19010 58212 19022
rect 58156 18958 58158 19010
rect 58210 18958 58212 19010
rect 58156 18900 58212 18958
rect 58156 18834 58212 18844
rect 57932 18228 57988 18238
rect 57932 17890 57988 18172
rect 57932 17838 57934 17890
rect 57986 17838 57988 17890
rect 57932 17826 57988 17838
rect 53004 17602 53060 17612
rect 55580 17668 55636 17678
rect 55580 17574 55636 17612
rect 51660 17502 51662 17554
rect 51714 17502 51716 17554
rect 51100 16830 51102 16882
rect 51154 16830 51156 16882
rect 51100 16818 51156 16830
rect 51212 17442 51268 17454
rect 51212 17390 51214 17442
rect 51266 17390 51268 17442
rect 50316 16770 50372 16782
rect 50316 16718 50318 16770
rect 50370 16718 50372 16770
rect 46844 16660 46900 16670
rect 46844 16566 46900 16604
rect 47628 16660 47684 16670
rect 46844 15540 46900 15550
rect 46844 15538 47348 15540
rect 46844 15486 46846 15538
rect 46898 15486 47348 15538
rect 46844 15484 47348 15486
rect 46844 15474 46900 15484
rect 46732 15426 46788 15438
rect 46732 15374 46734 15426
rect 46786 15374 46788 15426
rect 46508 15314 46564 15326
rect 46508 15262 46510 15314
rect 46562 15262 46564 15314
rect 46396 14644 46452 14654
rect 46396 13748 46452 14588
rect 46508 13972 46564 15262
rect 46508 13906 46564 13916
rect 46620 14868 46676 14878
rect 46396 13654 46452 13692
rect 45276 13356 45444 13412
rect 44492 12180 44548 12190
rect 44492 12086 44548 12124
rect 44044 10892 44324 10948
rect 45388 11506 45444 13356
rect 45388 11454 45390 11506
rect 45442 11454 45444 11506
rect 44044 10052 44100 10892
rect 45388 10052 45444 11454
rect 45948 13356 46340 13412
rect 44044 9996 44548 10052
rect 44044 9826 44100 9996
rect 44044 9774 44046 9826
rect 44098 9774 44100 9826
rect 44044 9762 44100 9774
rect 44156 9828 44212 9838
rect 44156 9734 44212 9772
rect 44268 9602 44324 9614
rect 44268 9550 44270 9602
rect 44322 9550 44324 9602
rect 44268 8820 44324 9550
rect 44492 9042 44548 9996
rect 45388 9986 45444 9996
rect 45836 11172 45892 11182
rect 45948 11172 46004 13356
rect 46620 12852 46676 14812
rect 46732 13860 46788 15374
rect 47292 15426 47348 15484
rect 47628 15428 47684 16604
rect 50204 16212 50260 16222
rect 50092 16100 50148 16110
rect 50092 15988 50148 16044
rect 50204 16098 50260 16156
rect 50204 16046 50206 16098
rect 50258 16046 50260 16098
rect 50204 16034 50260 16046
rect 49980 15986 50148 15988
rect 49980 15934 50094 15986
rect 50146 15934 50148 15986
rect 49980 15932 50148 15934
rect 49868 15876 49924 15886
rect 49868 15782 49924 15820
rect 47292 15374 47294 15426
rect 47346 15374 47348 15426
rect 47292 15362 47348 15374
rect 47516 15426 47684 15428
rect 47516 15374 47630 15426
rect 47682 15374 47684 15426
rect 47516 15372 47684 15374
rect 47068 15316 47124 15326
rect 47068 15222 47124 15260
rect 47068 14642 47124 14654
rect 47068 14590 47070 14642
rect 47122 14590 47124 14642
rect 47068 14308 47124 14590
rect 47516 14418 47572 15372
rect 47628 15362 47684 15372
rect 48300 15428 48356 15438
rect 48300 15334 48356 15372
rect 49868 14756 49924 14766
rect 49980 14756 50036 15932
rect 50092 15922 50148 15932
rect 49868 14754 50036 14756
rect 49868 14702 49870 14754
rect 49922 14702 50036 14754
rect 49868 14700 50036 14702
rect 48524 14532 48580 14542
rect 47516 14366 47518 14418
rect 47570 14366 47572 14418
rect 47516 14354 47572 14366
rect 47740 14530 48580 14532
rect 47740 14478 48526 14530
rect 48578 14478 48580 14530
rect 47740 14476 48580 14478
rect 47068 14242 47124 14252
rect 47404 13972 47460 13982
rect 47404 13878 47460 13916
rect 47628 13972 47684 13982
rect 47740 13972 47796 14476
rect 48524 14466 48580 14476
rect 47628 13970 47796 13972
rect 47628 13918 47630 13970
rect 47682 13918 47796 13970
rect 47628 13916 47796 13918
rect 47628 13906 47684 13916
rect 46732 13766 46788 13804
rect 47292 13748 47348 13786
rect 47292 13682 47348 13692
rect 49532 13748 49588 13758
rect 46844 13634 46900 13646
rect 46844 13582 46846 13634
rect 46898 13582 46900 13634
rect 46844 13076 46900 13582
rect 46844 13010 46900 13020
rect 47292 13524 47348 13534
rect 46620 12796 46788 12852
rect 46620 12178 46676 12190
rect 46620 12126 46622 12178
rect 46674 12126 46676 12178
rect 46620 12068 46676 12126
rect 46396 12012 46620 12068
rect 46396 11506 46452 12012
rect 46620 12002 46676 12012
rect 46732 12066 46788 12796
rect 46732 12014 46734 12066
rect 46786 12014 46788 12066
rect 46620 11620 46676 11630
rect 46732 11620 46788 12014
rect 46620 11618 46788 11620
rect 46620 11566 46622 11618
rect 46674 11566 46788 11618
rect 46620 11564 46788 11566
rect 46620 11554 46676 11564
rect 46396 11454 46398 11506
rect 46450 11454 46452 11506
rect 46396 11442 46452 11454
rect 46956 11506 47012 11518
rect 46956 11454 46958 11506
rect 47010 11454 47012 11506
rect 46956 11396 47012 11454
rect 46956 11330 47012 11340
rect 47292 11394 47348 13468
rect 49532 13186 49588 13692
rect 49868 13746 49924 14700
rect 49868 13694 49870 13746
rect 49922 13694 49924 13746
rect 49868 13682 49924 13694
rect 50316 13746 50372 16718
rect 51212 16212 51268 17390
rect 51660 16884 51716 17502
rect 58156 16994 58212 17006
rect 58156 16942 58158 16994
rect 58210 16942 58212 16994
rect 51772 16884 51828 16894
rect 51660 16882 51828 16884
rect 51660 16830 51774 16882
rect 51826 16830 51828 16882
rect 51660 16828 51828 16830
rect 51772 16818 51828 16828
rect 51884 16884 51940 16894
rect 51884 16660 51940 16828
rect 53116 16884 53172 16894
rect 53116 16790 53172 16828
rect 51212 16118 51268 16156
rect 51772 16604 51940 16660
rect 57932 16772 57988 16782
rect 50876 16100 50932 16110
rect 50876 16006 50932 16044
rect 51548 15988 51604 15998
rect 51548 15894 51604 15932
rect 50988 15876 51044 15886
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 50988 15426 51044 15820
rect 50988 15374 50990 15426
rect 51042 15374 51044 15426
rect 50988 15362 51044 15374
rect 51100 15428 51156 15438
rect 51100 15334 51156 15372
rect 51324 15314 51380 15326
rect 51324 15262 51326 15314
rect 51378 15262 51380 15314
rect 51324 15204 51380 15262
rect 51324 15138 51380 15148
rect 51772 15314 51828 16604
rect 57932 16322 57988 16716
rect 57932 16270 57934 16322
rect 57986 16270 57988 16322
rect 57932 16258 57988 16270
rect 58156 16212 58212 16942
rect 58156 16146 58212 16156
rect 53004 16100 53060 16110
rect 52668 15988 52724 15998
rect 52668 15894 52724 15932
rect 53004 15986 53060 16044
rect 55580 16100 55636 16110
rect 55580 16006 55636 16044
rect 53004 15934 53006 15986
rect 53058 15934 53060 15986
rect 53004 15922 53060 15934
rect 57932 15540 57988 15550
rect 51772 15262 51774 15314
rect 51826 15262 51828 15314
rect 51772 14980 51828 15262
rect 52332 15428 52388 15438
rect 51884 15204 51940 15214
rect 51884 15110 51940 15148
rect 51212 14924 51828 14980
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 50316 13694 50318 13746
rect 50370 13694 50372 13746
rect 50316 13682 50372 13694
rect 49532 13134 49534 13186
rect 49586 13134 49588 13186
rect 49532 13122 49588 13134
rect 50428 13634 50484 13646
rect 50428 13582 50430 13634
rect 50482 13582 50484 13634
rect 48972 13076 49028 13086
rect 48972 12982 49028 13020
rect 50092 13076 50148 13086
rect 49196 12964 49252 12974
rect 47516 12292 47572 12302
rect 47516 12198 47572 12236
rect 49196 12292 49252 12908
rect 49196 12226 49252 12236
rect 50092 12962 50148 13020
rect 50092 12910 50094 12962
rect 50146 12910 50148 12962
rect 50092 12178 50148 12910
rect 50092 12126 50094 12178
rect 50146 12126 50148 12178
rect 50092 12114 50148 12126
rect 50204 13074 50260 13086
rect 50204 13022 50206 13074
rect 50258 13022 50260 13074
rect 50204 12964 50260 13022
rect 50204 12180 50260 12908
rect 50316 12180 50372 12190
rect 50204 12178 50372 12180
rect 50204 12126 50318 12178
rect 50370 12126 50372 12178
rect 50204 12124 50372 12126
rect 50316 12114 50372 12124
rect 50428 11620 50484 13582
rect 50764 13188 50820 13198
rect 51212 13188 51268 14924
rect 51772 13972 51828 13982
rect 51324 13970 51828 13972
rect 51324 13918 51774 13970
rect 51826 13918 51828 13970
rect 51324 13916 51828 13918
rect 51324 13746 51380 13916
rect 51772 13906 51828 13916
rect 52332 13858 52388 15372
rect 53340 15426 53396 15438
rect 53340 15374 53342 15426
rect 53394 15374 53396 15426
rect 52668 15316 52724 15326
rect 53004 15316 53060 15326
rect 52668 15314 53060 15316
rect 52668 15262 52670 15314
rect 52722 15262 53006 15314
rect 53058 15262 53060 15314
rect 52668 15260 53060 15262
rect 52668 15250 52724 15260
rect 53004 15250 53060 15260
rect 53340 14532 53396 15374
rect 57932 14754 57988 15484
rect 57932 14702 57934 14754
rect 57986 14702 57988 14754
rect 57932 14690 57988 14702
rect 53340 14466 53396 14476
rect 55580 14532 55636 14542
rect 55580 14438 55636 14476
rect 52332 13806 52334 13858
rect 52386 13806 52388 13858
rect 52332 13794 52388 13806
rect 58156 13858 58212 13870
rect 58156 13806 58158 13858
rect 58210 13806 58212 13858
rect 51660 13748 51716 13758
rect 51324 13694 51326 13746
rect 51378 13694 51380 13746
rect 51324 13682 51380 13694
rect 51436 13746 51716 13748
rect 51436 13694 51662 13746
rect 51714 13694 51716 13746
rect 51436 13692 51716 13694
rect 50764 13186 51268 13188
rect 50764 13134 50766 13186
rect 50818 13134 51268 13186
rect 50764 13132 51268 13134
rect 50764 13122 50820 13132
rect 51436 13076 51492 13692
rect 51660 13682 51716 13692
rect 52220 13748 52276 13758
rect 52220 13654 52276 13692
rect 58156 13524 58212 13806
rect 58156 13458 58212 13468
rect 50876 13020 51492 13076
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 50652 12404 50708 12414
rect 50876 12404 50932 13020
rect 50652 12402 50932 12404
rect 50652 12350 50654 12402
rect 50706 12350 50932 12402
rect 50652 12348 50932 12350
rect 58156 12738 58212 12750
rect 58156 12686 58158 12738
rect 58210 12686 58212 12738
rect 50652 12338 50708 12348
rect 58156 12180 58212 12686
rect 58156 12114 58212 12124
rect 50204 11564 50484 11620
rect 50204 11506 50260 11564
rect 50204 11454 50206 11506
rect 50258 11454 50260 11506
rect 50204 11442 50260 11454
rect 47292 11342 47294 11394
rect 47346 11342 47348 11394
rect 47292 11330 47348 11342
rect 47516 11396 47572 11406
rect 47516 11302 47572 11340
rect 50316 11394 50372 11406
rect 50316 11342 50318 11394
rect 50370 11342 50372 11394
rect 45836 11170 46004 11172
rect 45836 11118 45838 11170
rect 45890 11118 46004 11170
rect 45836 11116 46004 11118
rect 47852 11172 47908 11182
rect 45052 9828 45108 9838
rect 45052 9734 45108 9772
rect 45388 9828 45444 9838
rect 45388 9714 45444 9772
rect 45388 9662 45390 9714
rect 45442 9662 45444 9714
rect 45388 9266 45444 9662
rect 45836 9714 45892 11116
rect 47852 11078 47908 11116
rect 48972 11172 49028 11182
rect 46732 10612 46788 10622
rect 46732 10518 46788 10556
rect 47180 10612 47236 10622
rect 47068 10498 47124 10510
rect 47068 10446 47070 10498
rect 47122 10446 47124 10498
rect 46284 9940 46340 9950
rect 46284 9846 46340 9884
rect 47068 9940 47124 10446
rect 47068 9846 47124 9884
rect 46508 9828 46564 9838
rect 46508 9734 46564 9772
rect 47180 9826 47236 10556
rect 47628 10612 47684 10622
rect 47628 10518 47684 10556
rect 48860 10612 48916 10622
rect 48860 10052 48916 10556
rect 48972 10612 49028 11116
rect 48972 10610 49252 10612
rect 48972 10558 48974 10610
rect 49026 10558 49252 10610
rect 48972 10556 49252 10558
rect 48972 10546 49028 10556
rect 48972 10052 49028 10062
rect 48860 10050 49028 10052
rect 48860 9998 48974 10050
rect 49026 9998 49028 10050
rect 48860 9996 49028 9998
rect 48972 9986 49028 9996
rect 47180 9774 47182 9826
rect 47234 9774 47236 9826
rect 47180 9762 47236 9774
rect 45836 9662 45838 9714
rect 45890 9662 45892 9714
rect 45836 9650 45892 9662
rect 47852 9714 47908 9726
rect 47852 9662 47854 9714
rect 47906 9662 47908 9714
rect 45388 9214 45390 9266
rect 45442 9214 45444 9266
rect 45388 9202 45444 9214
rect 47852 9156 47908 9662
rect 49196 9714 49252 10556
rect 49196 9662 49198 9714
rect 49250 9662 49252 9714
rect 49196 9650 49252 9662
rect 50204 10388 50260 10398
rect 50316 10388 50372 11342
rect 50204 10386 50372 10388
rect 50204 10334 50206 10386
rect 50258 10334 50372 10386
rect 50204 10332 50372 10334
rect 49084 9604 49140 9614
rect 49084 9510 49140 9548
rect 49980 9604 50036 9614
rect 44492 8990 44494 9042
rect 44546 8990 44548 9042
rect 44492 8978 44548 8990
rect 44940 9044 44996 9054
rect 44940 8950 44996 8988
rect 45612 9042 45668 9054
rect 45612 8990 45614 9042
rect 45666 8990 45668 9042
rect 44268 8754 44324 8764
rect 44716 8820 44772 8830
rect 44716 8726 44772 8764
rect 45612 8428 45668 8990
rect 43036 8194 43092 8204
rect 42700 8146 42980 8148
rect 42700 8094 42702 8146
rect 42754 8094 42980 8146
rect 42700 8092 42980 8094
rect 42700 7812 42756 8092
rect 42700 7746 42756 7756
rect 43372 8036 43428 8046
rect 42028 7634 42084 7644
rect 42252 7476 42308 7486
rect 42252 7382 42308 7420
rect 42812 7474 42868 7486
rect 42812 7422 42814 7474
rect 42866 7422 42868 7474
rect 41468 6290 41524 6300
rect 42140 7362 42196 7374
rect 42140 7310 42142 7362
rect 42194 7310 42196 7362
rect 41356 6132 41412 6142
rect 42140 6132 42196 7310
rect 42252 6132 42308 6142
rect 41356 6130 41636 6132
rect 41356 6078 41358 6130
rect 41410 6078 41636 6130
rect 41356 6076 41636 6078
rect 42140 6130 42308 6132
rect 42140 6078 42254 6130
rect 42306 6078 42308 6130
rect 42140 6076 42308 6078
rect 41356 6066 41412 6076
rect 41244 5908 41300 5918
rect 41244 5814 41300 5852
rect 41468 5906 41524 5918
rect 41468 5854 41470 5906
rect 41522 5854 41524 5906
rect 41468 5572 41524 5854
rect 41468 5506 41524 5516
rect 41580 5908 41636 6076
rect 42252 6066 42308 6076
rect 42812 6132 42868 7422
rect 43372 7474 43428 7980
rect 43372 7422 43374 7474
rect 43426 7422 43428 7474
rect 43372 7410 43428 7422
rect 43932 7474 43988 8316
rect 45388 8372 45444 8382
rect 45164 8260 45220 8270
rect 45164 8166 45220 8204
rect 45388 8258 45444 8316
rect 45388 8206 45390 8258
rect 45442 8206 45444 8258
rect 45388 8194 45444 8206
rect 45500 8372 45668 8428
rect 45836 9042 45892 9054
rect 45836 8990 45838 9042
rect 45890 8990 45892 9042
rect 45836 8482 45892 8990
rect 46172 9042 46228 9054
rect 46172 8990 46174 9042
rect 46226 8990 46228 9042
rect 45836 8430 45838 8482
rect 45890 8430 45892 8482
rect 45500 8370 45556 8372
rect 45500 8318 45502 8370
rect 45554 8318 45556 8370
rect 45500 8260 45556 8318
rect 45500 8194 45556 8204
rect 43932 7422 43934 7474
rect 43986 7422 43988 7474
rect 43932 7410 43988 7422
rect 45500 7924 45556 7934
rect 45500 7474 45556 7868
rect 45500 7422 45502 7474
rect 45554 7422 45556 7474
rect 45500 7410 45556 7422
rect 45836 7474 45892 8430
rect 45836 7422 45838 7474
rect 45890 7422 45892 7474
rect 45836 7410 45892 7422
rect 46060 8930 46116 8942
rect 46060 8878 46062 8930
rect 46114 8878 46116 8930
rect 43596 7250 43652 7262
rect 43596 7198 43598 7250
rect 43650 7198 43652 7250
rect 42812 6066 42868 6076
rect 43036 6076 43428 6132
rect 41692 5908 41748 5918
rect 41580 5906 41748 5908
rect 41580 5854 41694 5906
rect 41746 5854 41748 5906
rect 41580 5852 41748 5854
rect 41580 5290 41636 5852
rect 41692 5842 41748 5852
rect 42140 5906 42196 5918
rect 42140 5854 42142 5906
rect 42194 5854 42196 5906
rect 42140 5684 42196 5854
rect 41580 5238 41582 5290
rect 41634 5238 41636 5290
rect 41580 5226 41636 5238
rect 41916 5572 41972 5582
rect 41244 5124 41300 5134
rect 41244 5122 41412 5124
rect 41244 5070 41246 5122
rect 41298 5070 41412 5122
rect 41244 5068 41412 5070
rect 41244 5058 41300 5068
rect 41356 5012 41412 5068
rect 41804 5122 41860 5134
rect 41804 5070 41806 5122
rect 41858 5070 41860 5122
rect 41804 5012 41860 5070
rect 41356 4956 41860 5012
rect 41916 4900 41972 5516
rect 42140 5236 42196 5628
rect 42364 5906 42420 5918
rect 42364 5854 42366 5906
rect 42418 5854 42420 5906
rect 42364 5460 42420 5854
rect 42924 5684 42980 5694
rect 42924 5590 42980 5628
rect 42364 5394 42420 5404
rect 43036 5348 43092 6076
rect 43148 5908 43204 5918
rect 43372 5908 43428 6076
rect 43484 5908 43540 5918
rect 43372 5906 43540 5908
rect 43372 5854 43486 5906
rect 43538 5854 43540 5906
rect 43372 5852 43540 5854
rect 43148 5814 43204 5852
rect 43484 5842 43540 5852
rect 42140 5170 42196 5180
rect 42924 5292 43092 5348
rect 43260 5794 43316 5806
rect 43260 5742 43262 5794
rect 43314 5742 43316 5794
rect 42140 5012 42196 5022
rect 42140 4918 42196 4956
rect 41916 4834 41972 4844
rect 42924 4562 42980 5292
rect 43260 5234 43316 5742
rect 43596 5460 43652 7198
rect 44268 6132 44324 6142
rect 44268 6038 44324 6076
rect 44156 5906 44212 5918
rect 44156 5854 44158 5906
rect 44210 5854 44212 5906
rect 43708 5684 43764 5694
rect 43708 5590 43764 5628
rect 43596 5404 43876 5460
rect 43260 5182 43262 5234
rect 43314 5182 43316 5234
rect 43260 5170 43316 5182
rect 43036 5122 43092 5134
rect 43036 5070 43038 5122
rect 43090 5070 43092 5122
rect 43036 5012 43092 5070
rect 43708 5012 43764 5022
rect 43036 4946 43092 4956
rect 43372 5010 43764 5012
rect 43372 4958 43710 5010
rect 43762 4958 43764 5010
rect 43372 4956 43764 4958
rect 42924 4510 42926 4562
rect 42978 4510 42980 4562
rect 42924 4498 42980 4510
rect 42812 4452 42868 4462
rect 42812 4358 42868 4396
rect 43372 4338 43428 4956
rect 43708 4946 43764 4956
rect 43820 4788 43876 5404
rect 44156 5346 44212 5854
rect 44604 5908 44660 5918
rect 44604 5814 44660 5852
rect 46060 5908 46116 8878
rect 46172 7924 46228 8990
rect 46172 7858 46228 7868
rect 47068 7364 47124 7374
rect 47068 7270 47124 7308
rect 47852 6690 47908 9100
rect 49084 9156 49140 9166
rect 48188 8932 48244 8942
rect 48188 8258 48244 8876
rect 49084 8428 49140 9100
rect 49420 9042 49476 9054
rect 49420 8990 49422 9042
rect 49474 8990 49476 9042
rect 49196 8932 49252 8942
rect 49196 8838 49252 8876
rect 49084 8372 49364 8428
rect 48188 8206 48190 8258
rect 48242 8206 48244 8258
rect 48188 8194 48244 8206
rect 48524 8316 49028 8372
rect 48524 8258 48580 8316
rect 48524 8206 48526 8258
rect 48578 8206 48580 8258
rect 48524 8194 48580 8206
rect 48636 8146 48692 8158
rect 48636 8094 48638 8146
rect 48690 8094 48692 8146
rect 48300 7364 48356 7374
rect 48300 6802 48356 7308
rect 48300 6750 48302 6802
rect 48354 6750 48356 6802
rect 48300 6738 48356 6750
rect 47852 6638 47854 6690
rect 47906 6638 47908 6690
rect 47852 6626 47908 6638
rect 48636 6020 48692 8094
rect 48972 7586 49028 8316
rect 48972 7534 48974 7586
rect 49026 7534 49028 7586
rect 48972 7522 49028 7534
rect 49084 7476 49140 7486
rect 49084 6690 49140 7420
rect 49308 7474 49364 8372
rect 49308 7422 49310 7474
rect 49362 7422 49364 7474
rect 49308 7410 49364 7422
rect 49420 7364 49476 8990
rect 49532 9044 49588 9054
rect 49532 8258 49588 8988
rect 49980 9042 50036 9548
rect 49980 8990 49982 9042
rect 50034 8990 50036 9042
rect 49980 8978 50036 8990
rect 50204 9044 50260 10332
rect 50428 9156 50484 11564
rect 57932 11508 57988 11518
rect 57932 11414 57988 11452
rect 51660 11396 51716 11406
rect 50988 11284 51044 11294
rect 51324 11284 51380 11294
rect 50988 11282 51380 11284
rect 50988 11230 50990 11282
rect 51042 11230 51326 11282
rect 51378 11230 51380 11282
rect 50988 11228 51380 11230
rect 50988 11218 51044 11228
rect 51324 11218 51380 11228
rect 51660 11282 51716 11340
rect 55580 11396 55636 11406
rect 55580 11302 55636 11340
rect 51660 11230 51662 11282
rect 51714 11230 51716 11282
rect 51660 11218 51716 11230
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 58156 10836 58212 10846
rect 57708 10722 57764 10734
rect 57708 10670 57710 10722
rect 57762 10670 57764 10722
rect 57708 10164 57764 10670
rect 58156 10498 58212 10780
rect 58156 10446 58158 10498
rect 58210 10446 58212 10498
rect 58156 10434 58212 10446
rect 57708 10098 57764 10108
rect 51436 9604 51492 9614
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 51436 9266 51492 9548
rect 58156 9602 58212 9614
rect 58156 9550 58158 9602
rect 58210 9550 58212 9602
rect 58156 9492 58212 9550
rect 58156 9426 58212 9436
rect 51436 9214 51438 9266
rect 51490 9214 51492 9266
rect 51436 9202 51492 9214
rect 50540 9156 50596 9166
rect 50428 9154 50596 9156
rect 50428 9102 50542 9154
rect 50594 9102 50596 9154
rect 50428 9100 50596 9102
rect 50204 8978 50260 8988
rect 50540 8370 50596 9100
rect 50764 9154 50820 9166
rect 50764 9102 50766 9154
rect 50818 9102 50820 9154
rect 50652 9044 50708 9054
rect 50764 9044 50820 9102
rect 50708 8988 50820 9044
rect 50652 8978 50708 8988
rect 51324 8930 51380 8942
rect 51324 8878 51326 8930
rect 51378 8878 51380 8930
rect 50876 8820 50932 8830
rect 51212 8820 51268 8830
rect 50876 8818 51268 8820
rect 50876 8766 50878 8818
rect 50930 8766 51214 8818
rect 51266 8766 51268 8818
rect 50876 8764 51268 8766
rect 50876 8754 50932 8764
rect 51212 8754 51268 8764
rect 51324 8428 51380 8878
rect 50540 8318 50542 8370
rect 50594 8318 50596 8370
rect 50540 8306 50596 8318
rect 51212 8372 51380 8428
rect 57932 8372 57988 8382
rect 49532 8206 49534 8258
rect 49586 8206 49588 8258
rect 49532 8194 49588 8206
rect 50876 8258 50932 8270
rect 50876 8206 50878 8258
rect 50930 8206 50932 8258
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 50876 7476 50932 8206
rect 50876 7382 50932 7420
rect 51212 7474 51268 8372
rect 57932 8278 57988 8316
rect 51996 8260 52052 8270
rect 51660 8148 51716 8158
rect 51324 8146 51716 8148
rect 51324 8094 51662 8146
rect 51714 8094 51716 8146
rect 51324 8092 51716 8094
rect 51324 7586 51380 8092
rect 51660 8082 51716 8092
rect 51996 8146 52052 8204
rect 55580 8260 55636 8270
rect 55580 8166 55636 8204
rect 51996 8094 51998 8146
rect 52050 8094 52052 8146
rect 51996 8082 52052 8094
rect 58156 8148 58212 8158
rect 58156 7698 58212 8092
rect 58156 7646 58158 7698
rect 58210 7646 58212 7698
rect 58156 7634 58212 7646
rect 51324 7534 51326 7586
rect 51378 7534 51380 7586
rect 51324 7522 51380 7534
rect 51212 7422 51214 7474
rect 51266 7422 51268 7474
rect 51212 7410 51268 7422
rect 49420 7270 49476 7308
rect 49084 6638 49086 6690
rect 49138 6638 49140 6690
rect 49084 6626 49140 6638
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 48748 6020 48804 6030
rect 48524 5964 48748 6020
rect 46060 5842 46116 5852
rect 46732 5908 46788 5918
rect 46732 5814 46788 5852
rect 47628 5908 47684 5918
rect 47628 5814 47684 5852
rect 48412 5908 48468 5918
rect 45164 5794 45220 5806
rect 45164 5742 45166 5794
rect 45218 5742 45220 5794
rect 44156 5294 44158 5346
rect 44210 5294 44212 5346
rect 44156 5282 44212 5294
rect 44380 5684 44436 5694
rect 44380 5236 44436 5628
rect 44380 5170 44436 5180
rect 45164 5124 45220 5742
rect 46396 5794 46452 5806
rect 46396 5742 46398 5794
rect 46450 5742 46452 5794
rect 45164 5058 45220 5068
rect 45276 5682 45332 5694
rect 45276 5630 45278 5682
rect 45330 5630 45332 5682
rect 44044 5012 44100 5022
rect 44044 4918 44100 4956
rect 44156 4900 44212 4910
rect 44156 4806 44212 4844
rect 43820 4732 44100 4788
rect 43372 4286 43374 4338
rect 43426 4286 43428 4338
rect 43372 4274 43428 4286
rect 43596 4450 43652 4462
rect 43596 4398 43598 4450
rect 43650 4398 43652 4450
rect 43596 4340 43652 4398
rect 43932 4340 43988 4350
rect 43596 4338 43988 4340
rect 43596 4286 43934 4338
rect 43986 4286 43988 4338
rect 43596 4284 43988 4286
rect 43932 4274 43988 4284
rect 43708 4116 43764 4126
rect 41132 3266 41188 3276
rect 42364 3668 42420 3678
rect 30492 1586 30548 1596
rect 42364 800 42420 3612
rect 43708 800 43764 4060
rect 44044 3554 44100 4732
rect 45276 4676 45332 5630
rect 46396 5572 46452 5742
rect 46396 5506 46452 5516
rect 46508 5796 46564 5806
rect 46396 5348 46452 5358
rect 45948 5346 46452 5348
rect 45948 5294 46398 5346
rect 46450 5294 46452 5346
rect 45948 5292 46452 5294
rect 45388 5122 45444 5134
rect 45388 5070 45390 5122
rect 45442 5070 45444 5122
rect 45388 4900 45444 5070
rect 45948 5122 46004 5292
rect 46396 5282 46452 5292
rect 45948 5070 45950 5122
rect 46002 5070 46004 5122
rect 45948 5058 46004 5070
rect 46060 5124 46116 5134
rect 46060 5030 46116 5068
rect 46508 5012 46564 5740
rect 47292 5796 47348 5806
rect 47292 5702 47348 5740
rect 47852 5682 47908 5694
rect 47852 5630 47854 5682
rect 47906 5630 47908 5682
rect 47852 5572 47908 5630
rect 48188 5684 48244 5694
rect 48188 5590 48244 5628
rect 47852 5506 47908 5516
rect 46732 5236 46788 5246
rect 46732 5142 46788 5180
rect 48076 5236 48132 5246
rect 48076 5142 48132 5180
rect 47068 5124 47124 5134
rect 47068 5030 47124 5068
rect 46508 5010 46900 5012
rect 46508 4958 46510 5010
rect 46562 4958 46900 5010
rect 46508 4956 46900 4958
rect 46508 4946 46564 4956
rect 45388 4834 45444 4844
rect 45276 4610 45332 4620
rect 46844 4562 46900 4956
rect 48412 5010 48468 5852
rect 48524 5122 48580 5964
rect 48748 5926 48804 5964
rect 48860 6018 48916 6030
rect 48860 5966 48862 6018
rect 48914 5966 48916 6018
rect 48860 5908 48916 5966
rect 48860 5842 48916 5852
rect 49420 6020 49476 6030
rect 49420 5906 49476 5964
rect 50988 6020 51044 6030
rect 50988 6018 51156 6020
rect 50988 5966 50990 6018
rect 51042 5966 51156 6018
rect 50988 5964 51156 5966
rect 50988 5954 51044 5964
rect 49420 5854 49422 5906
rect 49474 5854 49476 5906
rect 49420 5842 49476 5854
rect 49644 5908 49700 5918
rect 49644 5814 49700 5852
rect 50316 5908 50372 5918
rect 50652 5908 50708 5918
rect 50316 5906 50708 5908
rect 50316 5854 50318 5906
rect 50370 5854 50654 5906
rect 50706 5854 50708 5906
rect 50316 5852 50708 5854
rect 50316 5842 50372 5852
rect 50652 5842 50708 5852
rect 48860 5684 48916 5694
rect 50092 5684 50148 5694
rect 48860 5682 49028 5684
rect 48860 5630 48862 5682
rect 48914 5630 49028 5682
rect 48860 5628 49028 5630
rect 48860 5618 48916 5628
rect 48524 5070 48526 5122
rect 48578 5070 48580 5122
rect 48524 5058 48580 5070
rect 48412 4958 48414 5010
rect 48466 4958 48468 5010
rect 48412 4946 48468 4958
rect 48972 5012 49028 5628
rect 49084 5124 49140 5134
rect 49532 5124 49588 5134
rect 49084 5122 49588 5124
rect 49084 5070 49086 5122
rect 49138 5070 49534 5122
rect 49586 5070 49588 5122
rect 49084 5068 49588 5070
rect 49084 5058 49140 5068
rect 49532 5058 49588 5068
rect 50092 5124 50148 5628
rect 50092 5030 50148 5068
rect 48972 4946 49028 4956
rect 50428 5010 50484 5022
rect 50428 4958 50430 5010
rect 50482 4958 50484 5010
rect 47404 4900 47460 4910
rect 47404 4898 47572 4900
rect 47404 4846 47406 4898
rect 47458 4846 47572 4898
rect 47404 4844 47572 4846
rect 47404 4834 47460 4844
rect 46844 4510 46846 4562
rect 46898 4510 46900 4562
rect 46844 4498 46900 4510
rect 47404 4676 47460 4686
rect 47404 4338 47460 4620
rect 47404 4286 47406 4338
rect 47458 4286 47460 4338
rect 47404 4274 47460 4286
rect 44940 4116 44996 4126
rect 44940 4022 44996 4060
rect 47180 4114 47236 4126
rect 47180 4062 47182 4114
rect 47234 4062 47236 4114
rect 47180 4004 47236 4062
rect 47180 3938 47236 3948
rect 44604 3668 44660 3678
rect 44604 3574 44660 3612
rect 44044 3502 44046 3554
rect 44098 3502 44100 3554
rect 44044 3490 44100 3502
rect 47516 3554 47572 4844
rect 49420 4898 49476 4910
rect 49420 4846 49422 4898
rect 49474 4846 49476 4898
rect 49084 4676 49140 4686
rect 49084 4450 49140 4620
rect 49084 4398 49086 4450
rect 49138 4398 49140 4450
rect 49084 4386 49140 4398
rect 48860 4228 48916 4238
rect 49420 4228 49476 4846
rect 49644 4898 49700 4910
rect 49644 4846 49646 4898
rect 49698 4846 49700 4898
rect 49644 4676 49700 4846
rect 49644 4610 49700 4620
rect 50428 4564 50484 4958
rect 50764 4900 50820 4938
rect 50988 4900 51044 4910
rect 50764 4834 50820 4844
rect 50876 4898 51044 4900
rect 50876 4846 50990 4898
rect 51042 4846 51044 4898
rect 50876 4844 51044 4846
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 50652 4564 50708 4574
rect 50428 4562 50708 4564
rect 50428 4510 50654 4562
rect 50706 4510 50708 4562
rect 50428 4508 50708 4510
rect 50652 4498 50708 4508
rect 50764 4452 50820 4462
rect 50876 4452 50932 4844
rect 50988 4834 51044 4844
rect 50764 4450 50932 4452
rect 50764 4398 50766 4450
rect 50818 4398 50932 4450
rect 50764 4396 50932 4398
rect 50764 4386 50820 4396
rect 51100 4340 51156 5964
rect 51212 5124 51268 5134
rect 51212 5010 51268 5068
rect 51212 4958 51214 5010
rect 51266 4958 51268 5010
rect 51212 4946 51268 4958
rect 51324 5012 51380 5022
rect 51324 4918 51380 4956
rect 51436 4900 51492 4910
rect 51324 4340 51380 4350
rect 51100 4338 51380 4340
rect 51100 4286 51326 4338
rect 51378 4286 51380 4338
rect 51100 4284 51380 4286
rect 51324 4274 51380 4284
rect 48860 4226 49476 4228
rect 48860 4174 48862 4226
rect 48914 4174 49476 4226
rect 48860 4172 49476 4174
rect 48860 4004 48916 4172
rect 48860 3938 48916 3948
rect 51100 4116 51156 4126
rect 47516 3502 47518 3554
rect 47570 3502 47572 3554
rect 47516 3490 47572 3502
rect 50428 3668 50484 3678
rect 46396 3444 46452 3454
rect 46396 800 46452 3388
rect 48972 3444 49028 3454
rect 48972 3350 49028 3388
rect 50428 800 50484 3612
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 51100 800 51156 4060
rect 51436 3554 51492 4844
rect 52332 4116 52388 4126
rect 52332 4022 52388 4060
rect 52220 3668 52276 3678
rect 52220 3574 52276 3612
rect 51436 3502 51438 3554
rect 51490 3502 51492 3554
rect 51436 3490 51492 3502
rect 52444 3332 52500 3342
rect 52444 800 52500 3276
rect 54124 3332 54180 3342
rect 54124 3238 54180 3276
rect 4704 0 4816 800
rect 9408 0 9520 800
rect 28896 0 29008 800
rect 42336 0 42448 800
rect 43680 0 43792 800
rect 46368 0 46480 800
rect 50400 0 50512 800
rect 51072 0 51184 800
rect 52416 0 52528 800
<< via2 >>
rect 26684 57820 26740 57876
rect 15036 57708 15092 57764
rect 13804 56194 13860 56196
rect 13804 56142 13806 56194
rect 13806 56142 13858 56194
rect 13858 56142 13860 56194
rect 13804 56140 13860 56142
rect 12572 56028 12628 56084
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 4172 55020 4228 55076
rect 4732 55074 4788 55076
rect 4732 55022 4734 55074
rect 4734 55022 4786 55074
rect 4786 55022 4788 55074
rect 4732 55020 4788 55022
rect 12460 55074 12516 55076
rect 12460 55022 12462 55074
rect 12462 55022 12514 55074
rect 12514 55022 12516 55074
rect 12460 55020 12516 55022
rect 1932 54460 1988 54516
rect 12012 54684 12068 54740
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 6524 54124 6580 54180
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 1708 51100 1764 51156
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 8316 53452 8372 53508
rect 8764 52274 8820 52276
rect 8764 52222 8766 52274
rect 8766 52222 8818 52274
rect 8818 52222 8820 52274
rect 8764 52220 8820 52222
rect 8540 52108 8596 52164
rect 8204 51324 8260 51380
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 4284 48748 4340 48804
rect 4732 48802 4788 48804
rect 4732 48750 4734 48802
rect 4734 48750 4786 48802
rect 4786 48750 4788 48802
rect 4732 48748 4788 48750
rect 5628 48748 5684 48804
rect 1932 48412 1988 48468
rect 1932 48018 1988 48020
rect 1932 47966 1934 48018
rect 1934 47966 1986 48018
rect 1986 47966 1988 48018
rect 1932 47964 1988 47966
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 4284 47292 4340 47348
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 1708 42364 1764 42420
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 1708 41298 1764 41300
rect 1708 41246 1710 41298
rect 1710 41246 1762 41298
rect 1762 41246 1764 41298
rect 1708 41244 1764 41246
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 1708 39004 1764 39060
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4284 37212 4340 37268
rect 2156 37042 2212 37044
rect 2156 36990 2158 37042
rect 2158 36990 2210 37042
rect 2210 36990 2212 37042
rect 2156 36988 2212 36990
rect 1932 36594 1988 36596
rect 1932 36542 1934 36594
rect 1934 36542 1986 36594
rect 1986 36542 1988 36594
rect 1932 36540 1988 36542
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 1708 35644 1764 35700
rect 4284 35698 4340 35700
rect 4284 35646 4286 35698
rect 4286 35646 4338 35698
rect 4338 35646 4340 35698
rect 4284 35644 4340 35646
rect 5516 35532 5572 35588
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 1932 34972 1988 35028
rect 6300 45778 6356 45780
rect 6300 45726 6302 45778
rect 6302 45726 6354 45778
rect 6354 45726 6356 45778
rect 6300 45724 6356 45726
rect 6076 45612 6132 45668
rect 8316 49810 8372 49812
rect 8316 49758 8318 49810
rect 8318 49758 8370 49810
rect 8370 49758 8372 49810
rect 8316 49756 8372 49758
rect 7868 48748 7924 48804
rect 8092 48466 8148 48468
rect 8092 48414 8094 48466
rect 8094 48414 8146 48466
rect 8146 48414 8148 48466
rect 8092 48412 8148 48414
rect 7308 47346 7364 47348
rect 7308 47294 7310 47346
rect 7310 47294 7362 47346
rect 7362 47294 7364 47346
rect 7308 47292 7364 47294
rect 6972 46508 7028 46564
rect 7644 46396 7700 46452
rect 7196 45890 7252 45892
rect 7196 45838 7198 45890
rect 7198 45838 7250 45890
rect 7250 45838 7252 45890
rect 7196 45836 7252 45838
rect 6524 45612 6580 45668
rect 7644 45724 7700 45780
rect 7868 44994 7924 44996
rect 7868 44942 7870 44994
rect 7870 44942 7922 44994
rect 7922 44942 7924 44994
rect 7868 44940 7924 44942
rect 6636 43538 6692 43540
rect 6636 43486 6638 43538
rect 6638 43486 6690 43538
rect 6690 43486 6692 43538
rect 6636 43484 6692 43486
rect 7308 41692 7364 41748
rect 6636 41132 6692 41188
rect 7084 41186 7140 41188
rect 7084 41134 7086 41186
rect 7086 41134 7138 41186
rect 7138 41134 7140 41186
rect 7084 41132 7140 41134
rect 6860 40796 6916 40852
rect 6636 39618 6692 39620
rect 6636 39566 6638 39618
rect 6638 39566 6690 39618
rect 6690 39566 6692 39618
rect 6636 39564 6692 39566
rect 7868 44098 7924 44100
rect 7868 44046 7870 44098
rect 7870 44046 7922 44098
rect 7922 44046 7924 44098
rect 7868 44044 7924 44046
rect 7420 40796 7476 40852
rect 7532 40514 7588 40516
rect 7532 40462 7534 40514
rect 7534 40462 7586 40514
rect 7586 40462 7588 40514
rect 7532 40460 7588 40462
rect 7308 40012 7364 40068
rect 7308 39618 7364 39620
rect 7308 39566 7310 39618
rect 7310 39566 7362 39618
rect 7362 39566 7364 39618
rect 7308 39564 7364 39566
rect 7532 39394 7588 39396
rect 7532 39342 7534 39394
rect 7534 39342 7586 39394
rect 7586 39342 7588 39394
rect 7532 39340 7588 39342
rect 9324 52162 9380 52164
rect 9324 52110 9326 52162
rect 9326 52110 9378 52162
rect 9378 52110 9380 52162
rect 9324 52108 9380 52110
rect 11900 54402 11956 54404
rect 11900 54350 11902 54402
rect 11902 54350 11954 54402
rect 11954 54350 11956 54402
rect 11900 54348 11956 54350
rect 10668 53452 10724 53508
rect 9772 53228 9828 53284
rect 10892 53340 10948 53396
rect 11900 53340 11956 53396
rect 11340 52892 11396 52948
rect 11116 52386 11172 52388
rect 11116 52334 11118 52386
rect 11118 52334 11170 52386
rect 11170 52334 11172 52386
rect 11116 52332 11172 52334
rect 10780 52220 10836 52276
rect 10332 52108 10388 52164
rect 9996 51490 10052 51492
rect 9996 51438 9998 51490
rect 9998 51438 10050 51490
rect 10050 51438 10052 51490
rect 9996 51436 10052 51438
rect 9548 51324 9604 51380
rect 9548 50706 9604 50708
rect 9548 50654 9550 50706
rect 9550 50654 9602 50706
rect 9602 50654 9604 50706
rect 9548 50652 9604 50654
rect 8876 49810 8932 49812
rect 8876 49758 8878 49810
rect 8878 49758 8930 49810
rect 8930 49758 8932 49810
rect 8876 49756 8932 49758
rect 8764 48748 8820 48804
rect 10108 50428 10164 50484
rect 9548 49810 9604 49812
rect 9548 49758 9550 49810
rect 9550 49758 9602 49810
rect 9602 49758 9604 49810
rect 9548 49756 9604 49758
rect 8652 47234 8708 47236
rect 8652 47182 8654 47234
rect 8654 47182 8706 47234
rect 8706 47182 8708 47234
rect 8652 47180 8708 47182
rect 8540 46450 8596 46452
rect 8540 46398 8542 46450
rect 8542 46398 8594 46450
rect 8594 46398 8596 46450
rect 8540 46396 8596 46398
rect 8092 45500 8148 45556
rect 8876 47180 8932 47236
rect 11452 51660 11508 51716
rect 11116 51378 11172 51380
rect 11116 51326 11118 51378
rect 11118 51326 11170 51378
rect 11170 51326 11172 51378
rect 11116 51324 11172 51326
rect 10444 50428 10500 50484
rect 10444 49420 10500 49476
rect 9548 48748 9604 48804
rect 8876 46450 8932 46452
rect 8876 46398 8878 46450
rect 8878 46398 8930 46450
rect 8930 46398 8932 46450
rect 8876 46396 8932 46398
rect 8876 45890 8932 45892
rect 8876 45838 8878 45890
rect 8878 45838 8930 45890
rect 8930 45838 8932 45890
rect 8876 45836 8932 45838
rect 8764 45778 8820 45780
rect 8764 45726 8766 45778
rect 8766 45726 8818 45778
rect 8818 45726 8820 45778
rect 8764 45724 8820 45726
rect 8092 43762 8148 43764
rect 8092 43710 8094 43762
rect 8094 43710 8146 43762
rect 8146 43710 8148 43762
rect 8092 43708 8148 43710
rect 8204 43484 8260 43540
rect 8316 42642 8372 42644
rect 8316 42590 8318 42642
rect 8318 42590 8370 42642
rect 8370 42590 8372 42642
rect 8316 42588 8372 42590
rect 8204 41746 8260 41748
rect 8204 41694 8206 41746
rect 8206 41694 8258 41746
rect 8258 41694 8260 41746
rect 8204 41692 8260 41694
rect 7980 40796 8036 40852
rect 8092 40178 8148 40180
rect 8092 40126 8094 40178
rect 8094 40126 8146 40178
rect 8146 40126 8148 40178
rect 8092 40124 8148 40126
rect 8204 39564 8260 39620
rect 8092 39340 8148 39396
rect 7980 39228 8036 39284
rect 7868 39116 7924 39172
rect 9212 46620 9268 46676
rect 9436 45666 9492 45668
rect 9436 45614 9438 45666
rect 9438 45614 9490 45666
rect 9490 45614 9492 45666
rect 9436 45612 9492 45614
rect 9548 45388 9604 45444
rect 9660 46620 9716 46676
rect 9548 43538 9604 43540
rect 9548 43486 9550 43538
rect 9550 43486 9602 43538
rect 9602 43486 9604 43538
rect 9548 43484 9604 43486
rect 8540 42194 8596 42196
rect 8540 42142 8542 42194
rect 8542 42142 8594 42194
rect 8594 42142 8596 42194
rect 8540 42140 8596 42142
rect 8428 40012 8484 40068
rect 8428 39228 8484 39284
rect 8876 40684 8932 40740
rect 8988 40236 9044 40292
rect 9884 48524 9940 48580
rect 10556 49196 10612 49252
rect 10668 48300 10724 48356
rect 11116 49196 11172 49252
rect 11116 48802 11172 48804
rect 11116 48750 11118 48802
rect 11118 48750 11170 48802
rect 11170 48750 11172 48802
rect 11116 48748 11172 48750
rect 10892 48412 10948 48468
rect 12460 54572 12516 54628
rect 12124 52946 12180 52948
rect 12124 52894 12126 52946
rect 12126 52894 12178 52946
rect 12178 52894 12180 52946
rect 12124 52892 12180 52894
rect 12348 52668 12404 52724
rect 12908 55916 12964 55972
rect 12796 55692 12852 55748
rect 12348 52444 12404 52500
rect 14140 55970 14196 55972
rect 14140 55918 14142 55970
rect 14142 55918 14194 55970
rect 14194 55918 14196 55970
rect 14140 55916 14196 55918
rect 14140 55410 14196 55412
rect 14140 55358 14142 55410
rect 14142 55358 14194 55410
rect 14194 55358 14196 55410
rect 14140 55356 14196 55358
rect 25004 57484 25060 57540
rect 22988 57372 23044 57428
rect 21084 57260 21140 57316
rect 16380 57148 16436 57204
rect 15596 56140 15652 56196
rect 14588 55244 14644 55300
rect 14924 55244 14980 55300
rect 12908 54684 12964 54740
rect 14252 54460 14308 54516
rect 12908 54012 12964 54068
rect 13132 53900 13188 53956
rect 12572 52946 12628 52948
rect 12572 52894 12574 52946
rect 12574 52894 12626 52946
rect 12626 52894 12628 52946
rect 12572 52892 12628 52894
rect 12460 52332 12516 52388
rect 12348 51660 12404 51716
rect 12684 51378 12740 51380
rect 12684 51326 12686 51378
rect 12686 51326 12738 51378
rect 12738 51326 12740 51378
rect 12684 51324 12740 51326
rect 12236 50540 12292 50596
rect 11676 50092 11732 50148
rect 11452 49308 11508 49364
rect 11564 48972 11620 49028
rect 9996 47234 10052 47236
rect 9996 47182 9998 47234
rect 9998 47182 10050 47234
rect 10050 47182 10052 47234
rect 9996 47180 10052 47182
rect 9884 45836 9940 45892
rect 10332 46674 10388 46676
rect 10332 46622 10334 46674
rect 10334 46622 10386 46674
rect 10386 46622 10388 46674
rect 10332 46620 10388 46622
rect 9996 45052 10052 45108
rect 10444 45836 10500 45892
rect 10332 43932 10388 43988
rect 9772 41132 9828 41188
rect 10332 41916 10388 41972
rect 9660 40796 9716 40852
rect 9772 40908 9828 40964
rect 9212 40124 9268 40180
rect 9884 40626 9940 40628
rect 9884 40574 9886 40626
rect 9886 40574 9938 40626
rect 9938 40574 9940 40626
rect 9884 40572 9940 40574
rect 10220 40514 10276 40516
rect 10220 40462 10222 40514
rect 10222 40462 10274 40514
rect 10274 40462 10276 40514
rect 10220 40460 10276 40462
rect 10108 40402 10164 40404
rect 10108 40350 10110 40402
rect 10110 40350 10162 40402
rect 10162 40350 10164 40402
rect 10108 40348 10164 40350
rect 9996 39618 10052 39620
rect 9996 39566 9998 39618
rect 9998 39566 10050 39618
rect 10050 39566 10052 39618
rect 9996 39564 10052 39566
rect 9996 38892 10052 38948
rect 10332 39116 10388 39172
rect 8316 37884 8372 37940
rect 7196 37266 7252 37268
rect 7196 37214 7198 37266
rect 7198 37214 7250 37266
rect 7250 37214 7252 37266
rect 7196 37212 7252 37214
rect 8428 37212 8484 37268
rect 6412 36876 6468 36932
rect 8204 36428 8260 36484
rect 7420 36092 7476 36148
rect 6860 35532 6916 35588
rect 6300 34690 6356 34692
rect 6300 34638 6302 34690
rect 6302 34638 6354 34690
rect 6354 34638 6356 34690
rect 6300 34636 6356 34638
rect 5628 34412 5684 34468
rect 6076 34188 6132 34244
rect 4844 34076 4900 34132
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 2044 33234 2100 33236
rect 2044 33182 2046 33234
rect 2046 33182 2098 33234
rect 2098 33182 2100 33234
rect 2044 33180 2100 33182
rect 1708 32956 1764 33012
rect 2492 32956 2548 33012
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 2380 31666 2436 31668
rect 2380 31614 2382 31666
rect 2382 31614 2434 31666
rect 2434 31614 2436 31666
rect 2380 31612 2436 31614
rect 2044 31554 2100 31556
rect 2044 31502 2046 31554
rect 2046 31502 2098 31554
rect 2098 31502 2100 31554
rect 2044 31500 2100 31502
rect 1820 30940 1876 30996
rect 5516 34130 5572 34132
rect 5516 34078 5518 34130
rect 5518 34078 5570 34130
rect 5570 34078 5572 34130
rect 5516 34076 5572 34078
rect 6636 33852 6692 33908
rect 4284 30716 4340 30772
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 1932 30268 1988 30324
rect 2492 29596 2548 29652
rect 1932 29202 1988 29204
rect 1932 29150 1934 29202
rect 1934 29150 1986 29202
rect 1986 29150 1988 29202
rect 1932 29148 1988 29150
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4284 28812 4340 28868
rect 4284 28642 4340 28644
rect 4284 28590 4286 28642
rect 4286 28590 4338 28642
rect 4338 28590 4340 28642
rect 4284 28588 4340 28590
rect 4172 28476 4228 28532
rect 1932 28252 1988 28308
rect 7868 36258 7924 36260
rect 7868 36206 7870 36258
rect 7870 36206 7922 36258
rect 7922 36206 7924 36258
rect 7868 36204 7924 36206
rect 7532 33180 7588 33236
rect 7868 34636 7924 34692
rect 6636 30940 6692 30996
rect 8428 34748 8484 34804
rect 8540 35308 8596 35364
rect 8316 34636 8372 34692
rect 8316 34354 8372 34356
rect 8316 34302 8318 34354
rect 8318 34302 8370 34354
rect 8370 34302 8372 34354
rect 8316 34300 8372 34302
rect 8092 33964 8148 34020
rect 8316 34076 8372 34132
rect 10220 37938 10276 37940
rect 10220 37886 10222 37938
rect 10222 37886 10274 37938
rect 10274 37886 10276 37938
rect 10220 37884 10276 37886
rect 8988 36594 9044 36596
rect 8988 36542 8990 36594
rect 8990 36542 9042 36594
rect 9042 36542 9044 36594
rect 8988 36540 9044 36542
rect 8988 35644 9044 35700
rect 9436 35308 9492 35364
rect 9996 37212 10052 37268
rect 11452 47740 11508 47796
rect 11452 47570 11508 47572
rect 11452 47518 11454 47570
rect 11454 47518 11506 47570
rect 11506 47518 11508 47570
rect 11452 47516 11508 47518
rect 11452 47068 11508 47124
rect 11676 47628 11732 47684
rect 12012 49420 12068 49476
rect 12572 49196 12628 49252
rect 12236 48748 12292 48804
rect 11228 45276 11284 45332
rect 11228 43932 11284 43988
rect 10668 42700 10724 42756
rect 10668 41916 10724 41972
rect 10556 40908 10612 40964
rect 10668 40236 10724 40292
rect 10668 39676 10724 39732
rect 11116 41692 11172 41748
rect 11004 40908 11060 40964
rect 10892 40460 10948 40516
rect 10556 37826 10612 37828
rect 10556 37774 10558 37826
rect 10558 37774 10610 37826
rect 10610 37774 10612 37826
rect 10556 37772 10612 37774
rect 10444 37548 10500 37604
rect 10668 37266 10724 37268
rect 10668 37214 10670 37266
rect 10670 37214 10722 37266
rect 10722 37214 10724 37266
rect 10668 37212 10724 37214
rect 8764 34972 8820 35028
rect 8652 34914 8708 34916
rect 8652 34862 8654 34914
rect 8654 34862 8706 34914
rect 8706 34862 8708 34914
rect 8652 34860 8708 34862
rect 9436 34802 9492 34804
rect 9436 34750 9438 34802
rect 9438 34750 9490 34802
rect 9490 34750 9492 34802
rect 9436 34748 9492 34750
rect 8988 34636 9044 34692
rect 10444 36204 10500 36260
rect 10108 35644 10164 35700
rect 12012 46674 12068 46676
rect 12012 46622 12014 46674
rect 12014 46622 12066 46674
rect 12066 46622 12068 46674
rect 12012 46620 12068 46622
rect 11900 46508 11956 46564
rect 11564 46060 11620 46116
rect 11676 45836 11732 45892
rect 11788 45724 11844 45780
rect 11788 45276 11844 45332
rect 11788 44380 11844 44436
rect 11452 42140 11508 42196
rect 11564 42700 11620 42756
rect 11340 41970 11396 41972
rect 11340 41918 11342 41970
rect 11342 41918 11394 41970
rect 11394 41918 11396 41970
rect 11340 41916 11396 41918
rect 11340 41020 11396 41076
rect 11452 40348 11508 40404
rect 11676 42252 11732 42308
rect 11564 39340 11620 39396
rect 11676 40348 11732 40404
rect 11228 38668 11284 38724
rect 12348 48524 12404 48580
rect 12348 48188 12404 48244
rect 12460 48300 12516 48356
rect 12348 46508 12404 46564
rect 11900 43932 11956 43988
rect 13020 50204 13076 50260
rect 13580 54402 13636 54404
rect 13580 54350 13582 54402
rect 13582 54350 13634 54402
rect 13634 54350 13636 54402
rect 13580 54348 13636 54350
rect 13356 53564 13412 53620
rect 13692 53228 13748 53284
rect 13356 53170 13412 53172
rect 13356 53118 13358 53170
rect 13358 53118 13410 53170
rect 13410 53118 13412 53170
rect 13356 53116 13412 53118
rect 13244 51324 13300 51380
rect 13132 47404 13188 47460
rect 12908 45948 12964 46004
rect 13020 46956 13076 47012
rect 12684 44380 12740 44436
rect 13580 50764 13636 50820
rect 13916 52892 13972 52948
rect 13804 52834 13860 52836
rect 13804 52782 13806 52834
rect 13806 52782 13858 52834
rect 13858 52782 13860 52834
rect 13804 52780 13860 52782
rect 14252 52946 14308 52948
rect 14252 52894 14254 52946
rect 14254 52894 14306 52946
rect 14306 52894 14308 52946
rect 14252 52892 14308 52894
rect 13580 49196 13636 49252
rect 13692 50594 13748 50596
rect 13692 50542 13694 50594
rect 13694 50542 13746 50594
rect 13746 50542 13748 50594
rect 13692 50540 13748 50542
rect 13580 49026 13636 49028
rect 13580 48974 13582 49026
rect 13582 48974 13634 49026
rect 13634 48974 13636 49026
rect 13580 48972 13636 48974
rect 13468 48412 13524 48468
rect 13356 46956 13412 47012
rect 13580 46956 13636 47012
rect 13020 44940 13076 44996
rect 13356 45106 13412 45108
rect 13356 45054 13358 45106
rect 13358 45054 13410 45106
rect 13410 45054 13412 45106
rect 13356 45052 13412 45054
rect 12908 44322 12964 44324
rect 12908 44270 12910 44322
rect 12910 44270 12962 44322
rect 12962 44270 12964 44322
rect 12908 44268 12964 44270
rect 12124 41970 12180 41972
rect 12124 41918 12126 41970
rect 12126 41918 12178 41970
rect 12178 41918 12180 41970
rect 12124 41916 12180 41918
rect 12796 43820 12852 43876
rect 11900 39618 11956 39620
rect 11900 39566 11902 39618
rect 11902 39566 11954 39618
rect 11954 39566 11956 39618
rect 11900 39564 11956 39566
rect 11900 39004 11956 39060
rect 12684 42924 12740 42980
rect 12572 42812 12628 42868
rect 12460 41970 12516 41972
rect 12460 41918 12462 41970
rect 12462 41918 12514 41970
rect 12514 41918 12516 41970
rect 12460 41916 12516 41918
rect 12684 41804 12740 41860
rect 12684 41020 12740 41076
rect 12572 39058 12628 39060
rect 12572 39006 12574 39058
rect 12574 39006 12626 39058
rect 12626 39006 12628 39058
rect 12572 39004 12628 39006
rect 12236 38834 12292 38836
rect 12236 38782 12238 38834
rect 12238 38782 12290 38834
rect 12290 38782 12292 38834
rect 12236 38780 12292 38782
rect 12796 40236 12852 40292
rect 13580 44098 13636 44100
rect 13580 44046 13582 44098
rect 13582 44046 13634 44098
rect 13634 44046 13636 44098
rect 13580 44044 13636 44046
rect 14028 52108 14084 52164
rect 14476 54572 14532 54628
rect 15260 55356 15316 55412
rect 14700 54460 14756 54516
rect 14364 52220 14420 52276
rect 14476 53452 14532 53508
rect 14140 51324 14196 51380
rect 14812 53506 14868 53508
rect 14812 53454 14814 53506
rect 14814 53454 14866 53506
rect 14866 53454 14868 53506
rect 14812 53452 14868 53454
rect 14252 50652 14308 50708
rect 13804 49980 13860 50036
rect 13804 44882 13860 44884
rect 13804 44830 13806 44882
rect 13806 44830 13858 44882
rect 13858 44830 13860 44882
rect 13804 44828 13860 44830
rect 13804 44044 13860 44100
rect 14700 49196 14756 49252
rect 14028 46786 14084 46788
rect 14028 46734 14030 46786
rect 14030 46734 14082 46786
rect 14082 46734 14084 46786
rect 14028 46732 14084 46734
rect 14588 48972 14644 49028
rect 14476 48300 14532 48356
rect 14476 47292 14532 47348
rect 15372 55244 15428 55300
rect 15932 55298 15988 55300
rect 15932 55246 15934 55298
rect 15934 55246 15986 55298
rect 15986 55246 15988 55298
rect 15932 55244 15988 55246
rect 15596 55132 15652 55188
rect 15372 54572 15428 54628
rect 15260 51436 15316 51492
rect 14812 48076 14868 48132
rect 15036 50706 15092 50708
rect 15036 50654 15038 50706
rect 15038 50654 15090 50706
rect 15090 50654 15092 50706
rect 15036 50652 15092 50654
rect 15260 50034 15316 50036
rect 15260 49982 15262 50034
rect 15262 49982 15314 50034
rect 15314 49982 15316 50034
rect 15260 49980 15316 49982
rect 15260 49532 15316 49588
rect 15708 53730 15764 53732
rect 15708 53678 15710 53730
rect 15710 53678 15762 53730
rect 15762 53678 15764 53730
rect 15708 53676 15764 53678
rect 15484 53116 15540 53172
rect 15484 51996 15540 52052
rect 15484 51436 15540 51492
rect 16268 54402 16324 54404
rect 16268 54350 16270 54402
rect 16270 54350 16322 54402
rect 16322 54350 16324 54402
rect 16268 54348 16324 54350
rect 18284 56588 18340 56644
rect 18172 56252 18228 56308
rect 17836 56140 17892 56196
rect 16604 55244 16660 55300
rect 16492 55020 16548 55076
rect 16716 54572 16772 54628
rect 16492 53900 16548 53956
rect 16380 52834 16436 52836
rect 16380 52782 16382 52834
rect 16382 52782 16434 52834
rect 16434 52782 16436 52834
rect 16380 52780 16436 52782
rect 16044 52668 16100 52724
rect 16156 52162 16212 52164
rect 16156 52110 16158 52162
rect 16158 52110 16210 52162
rect 16210 52110 16212 52162
rect 16156 52108 16212 52110
rect 16156 51436 16212 51492
rect 15596 50594 15652 50596
rect 15596 50542 15598 50594
rect 15598 50542 15650 50594
rect 15650 50542 15652 50594
rect 15596 50540 15652 50542
rect 15708 49026 15764 49028
rect 15708 48974 15710 49026
rect 15710 48974 15762 49026
rect 15762 48974 15764 49026
rect 15708 48972 15764 48974
rect 15372 48412 15428 48468
rect 15820 48860 15876 48916
rect 15596 48242 15652 48244
rect 15596 48190 15598 48242
rect 15598 48190 15650 48242
rect 15650 48190 15652 48242
rect 15596 48188 15652 48190
rect 15820 47458 15876 47460
rect 15820 47406 15822 47458
rect 15822 47406 15874 47458
rect 15874 47406 15876 47458
rect 15820 47404 15876 47406
rect 15484 47068 15540 47124
rect 15260 46508 15316 46564
rect 14140 45724 14196 45780
rect 14140 45388 14196 45444
rect 14812 45388 14868 45444
rect 14812 44546 14868 44548
rect 14812 44494 14814 44546
rect 14814 44494 14866 44546
rect 14866 44494 14868 44546
rect 14812 44492 14868 44494
rect 14028 44268 14084 44324
rect 14028 44098 14084 44100
rect 14028 44046 14030 44098
rect 14030 44046 14082 44098
rect 14082 44046 14084 44098
rect 14028 44044 14084 44046
rect 13356 41804 13412 41860
rect 14476 44044 14532 44100
rect 14364 43650 14420 43652
rect 14364 43598 14366 43650
rect 14366 43598 14418 43650
rect 14418 43598 14420 43650
rect 14364 43596 14420 43598
rect 14140 43484 14196 43540
rect 14700 44098 14756 44100
rect 14700 44046 14702 44098
rect 14702 44046 14754 44098
rect 14754 44046 14756 44098
rect 14700 44044 14756 44046
rect 15148 44098 15204 44100
rect 15148 44046 15150 44098
rect 15150 44046 15202 44098
rect 15202 44046 15204 44098
rect 15148 44044 15204 44046
rect 14700 43708 14756 43764
rect 13804 41916 13860 41972
rect 14588 41970 14644 41972
rect 14588 41918 14590 41970
rect 14590 41918 14642 41970
rect 14642 41918 14644 41970
rect 14588 41916 14644 41918
rect 14924 43484 14980 43540
rect 14924 42140 14980 42196
rect 14924 41970 14980 41972
rect 14924 41918 14926 41970
rect 14926 41918 14978 41970
rect 14978 41918 14980 41970
rect 14924 41916 14980 41918
rect 15484 45948 15540 46004
rect 15484 44380 15540 44436
rect 16044 47852 16100 47908
rect 16380 51212 16436 51268
rect 16380 50428 16436 50484
rect 16268 49644 16324 49700
rect 16380 48860 16436 48916
rect 16156 47628 16212 47684
rect 16044 46956 16100 47012
rect 15932 46284 15988 46340
rect 15484 43932 15540 43988
rect 15708 44828 15764 44884
rect 15820 44604 15876 44660
rect 15708 44322 15764 44324
rect 15708 44270 15710 44322
rect 15710 44270 15762 44322
rect 15762 44270 15764 44322
rect 15708 44268 15764 44270
rect 15596 43484 15652 43540
rect 15260 42252 15316 42308
rect 14364 41186 14420 41188
rect 14364 41134 14366 41186
rect 14366 41134 14418 41186
rect 14418 41134 14420 41186
rect 14364 41132 14420 41134
rect 15148 41804 15204 41860
rect 14140 40348 14196 40404
rect 13468 39676 13524 39732
rect 13132 38722 13188 38724
rect 13132 38670 13134 38722
rect 13134 38670 13186 38722
rect 13186 38670 13188 38722
rect 13132 38668 13188 38670
rect 11788 36594 11844 36596
rect 11788 36542 11790 36594
rect 11790 36542 11842 36594
rect 11842 36542 11844 36594
rect 11788 36540 11844 36542
rect 12348 36482 12404 36484
rect 12348 36430 12350 36482
rect 12350 36430 12402 36482
rect 12402 36430 12404 36482
rect 12348 36428 12404 36430
rect 11116 36092 11172 36148
rect 13468 37826 13524 37828
rect 13468 37774 13470 37826
rect 13470 37774 13522 37826
rect 13522 37774 13524 37826
rect 13468 37772 13524 37774
rect 14028 39452 14084 39508
rect 14924 40572 14980 40628
rect 14700 40348 14756 40404
rect 14812 40124 14868 40180
rect 14924 39900 14980 39956
rect 14924 39676 14980 39732
rect 14812 39452 14868 39508
rect 14700 39228 14756 39284
rect 14364 38892 14420 38948
rect 14924 39116 14980 39172
rect 15148 40572 15204 40628
rect 15372 41244 15428 41300
rect 15708 42700 15764 42756
rect 16380 47180 16436 47236
rect 16268 46786 16324 46788
rect 16268 46734 16270 46786
rect 16270 46734 16322 46786
rect 16322 46734 16324 46786
rect 16268 46732 16324 46734
rect 17052 54236 17108 54292
rect 17052 54012 17108 54068
rect 16828 51100 16884 51156
rect 17164 53452 17220 53508
rect 17836 55916 17892 55972
rect 17388 55186 17444 55188
rect 17388 55134 17390 55186
rect 17390 55134 17442 55186
rect 17442 55134 17444 55186
rect 17388 55132 17444 55134
rect 17836 54460 17892 54516
rect 17388 54012 17444 54068
rect 17276 52780 17332 52836
rect 17052 52444 17108 52500
rect 16716 50876 16772 50932
rect 16940 50764 16996 50820
rect 17164 52556 17220 52612
rect 16604 50092 16660 50148
rect 16604 48748 16660 48804
rect 16828 50204 16884 50260
rect 16828 49868 16884 49924
rect 16828 48972 16884 49028
rect 16716 48636 16772 48692
rect 16828 48300 16884 48356
rect 16828 47404 16884 47460
rect 16492 46844 16548 46900
rect 16492 46562 16548 46564
rect 16492 46510 16494 46562
rect 16494 46510 16546 46562
rect 16546 46510 16548 46562
rect 16492 46508 16548 46510
rect 16828 46898 16884 46900
rect 16828 46846 16830 46898
rect 16830 46846 16882 46898
rect 16882 46846 16884 46898
rect 16828 46844 16884 46846
rect 16828 46172 16884 46228
rect 16380 44268 16436 44324
rect 15260 39004 15316 39060
rect 14252 38332 14308 38388
rect 16156 42588 16212 42644
rect 16268 44156 16324 44212
rect 16268 41468 16324 41524
rect 16380 43372 16436 43428
rect 16268 41132 16324 41188
rect 16716 45164 16772 45220
rect 16716 44492 16772 44548
rect 16828 44828 16884 44884
rect 18060 55522 18116 55524
rect 18060 55470 18062 55522
rect 18062 55470 18114 55522
rect 18114 55470 18116 55522
rect 18060 55468 18116 55470
rect 19628 56588 19684 56644
rect 19180 56194 19236 56196
rect 19180 56142 19182 56194
rect 19182 56142 19234 56194
rect 19234 56142 19236 56194
rect 19180 56140 19236 56142
rect 18844 55970 18900 55972
rect 18844 55918 18846 55970
rect 18846 55918 18898 55970
rect 18898 55918 18900 55970
rect 18844 55916 18900 55918
rect 18844 55692 18900 55748
rect 18732 55298 18788 55300
rect 18732 55246 18734 55298
rect 18734 55246 18786 55298
rect 18786 55246 18788 55298
rect 18732 55244 18788 55246
rect 18396 54460 18452 54516
rect 19180 55858 19236 55860
rect 19180 55806 19182 55858
rect 19182 55806 19234 55858
rect 19234 55806 19236 55858
rect 19180 55804 19236 55806
rect 19068 55522 19124 55524
rect 19068 55470 19070 55522
rect 19070 55470 19122 55522
rect 19122 55470 19124 55522
rect 19068 55468 19124 55470
rect 19180 55580 19236 55636
rect 18172 54236 18228 54292
rect 18060 53842 18116 53844
rect 18060 53790 18062 53842
rect 18062 53790 18114 53842
rect 18114 53790 18116 53842
rect 18060 53788 18116 53790
rect 17500 53340 17556 53396
rect 17500 53170 17556 53172
rect 17500 53118 17502 53170
rect 17502 53118 17554 53170
rect 17554 53118 17556 53170
rect 17500 53116 17556 53118
rect 17836 53228 17892 53284
rect 17612 52274 17668 52276
rect 17612 52222 17614 52274
rect 17614 52222 17666 52274
rect 17666 52222 17668 52274
rect 17612 52220 17668 52222
rect 17724 51378 17780 51380
rect 17724 51326 17726 51378
rect 17726 51326 17778 51378
rect 17778 51326 17780 51378
rect 17724 51324 17780 51326
rect 17500 50594 17556 50596
rect 17500 50542 17502 50594
rect 17502 50542 17554 50594
rect 17554 50542 17556 50594
rect 17500 50540 17556 50542
rect 18060 52332 18116 52388
rect 18844 53452 18900 53508
rect 18620 52668 18676 52724
rect 18284 52556 18340 52612
rect 18284 51996 18340 52052
rect 18060 51884 18116 51940
rect 18060 51436 18116 51492
rect 17948 51324 18004 51380
rect 19180 52220 19236 52276
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 20972 56140 21028 56196
rect 20188 56028 20244 56084
rect 19740 55468 19796 55524
rect 20188 55244 20244 55300
rect 20412 56028 20468 56084
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 19740 54514 19796 54516
rect 19740 54462 19742 54514
rect 19742 54462 19794 54514
rect 19794 54462 19796 54514
rect 19740 54460 19796 54462
rect 19628 54012 19684 54068
rect 19404 53954 19460 53956
rect 19404 53902 19406 53954
rect 19406 53902 19458 53954
rect 19458 53902 19460 53954
rect 19404 53900 19460 53902
rect 19404 53004 19460 53060
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 19740 52780 19796 52836
rect 20188 52780 20244 52836
rect 20748 55356 20804 55412
rect 20412 53842 20468 53844
rect 20412 53790 20414 53842
rect 20414 53790 20466 53842
rect 20466 53790 20468 53842
rect 20412 53788 20468 53790
rect 19628 52220 19684 52276
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 18732 51548 18788 51604
rect 19180 51378 19236 51380
rect 19180 51326 19182 51378
rect 19182 51326 19234 51378
rect 19234 51326 19236 51378
rect 19180 51324 19236 51326
rect 18844 51212 18900 51268
rect 18060 50540 18116 50596
rect 17388 49980 17444 50036
rect 17276 48300 17332 48356
rect 17388 49810 17444 49812
rect 17388 49758 17390 49810
rect 17390 49758 17442 49810
rect 17442 49758 17444 49810
rect 17388 49756 17444 49758
rect 17500 49026 17556 49028
rect 17500 48974 17502 49026
rect 17502 48974 17554 49026
rect 17554 48974 17556 49026
rect 17500 48972 17556 48974
rect 17052 47570 17108 47572
rect 17052 47518 17054 47570
rect 17054 47518 17106 47570
rect 17106 47518 17108 47570
rect 17052 47516 17108 47518
rect 17052 46620 17108 46676
rect 16828 44156 16884 44212
rect 16940 40684 16996 40740
rect 17388 47404 17444 47460
rect 17724 48914 17780 48916
rect 17724 48862 17726 48914
rect 17726 48862 17778 48914
rect 17778 48862 17780 48914
rect 17724 48860 17780 48862
rect 17612 46620 17668 46676
rect 17724 48636 17780 48692
rect 17724 47404 17780 47460
rect 17276 44156 17332 44212
rect 17500 45500 17556 45556
rect 18620 50540 18676 50596
rect 18732 51100 18788 51156
rect 18732 50652 18788 50708
rect 18284 49698 18340 49700
rect 18284 49646 18286 49698
rect 18286 49646 18338 49698
rect 18338 49646 18340 49698
rect 18284 49644 18340 49646
rect 17948 47852 18004 47908
rect 18284 47740 18340 47796
rect 18060 47068 18116 47124
rect 18284 47292 18340 47348
rect 18172 46956 18228 47012
rect 17836 46172 17892 46228
rect 17724 44604 17780 44660
rect 17052 42588 17108 42644
rect 16492 40626 16548 40628
rect 16492 40574 16494 40626
rect 16494 40574 16546 40626
rect 16546 40574 16548 40626
rect 16492 40572 16548 40574
rect 16268 40348 16324 40404
rect 15820 40236 15876 40292
rect 16940 40236 16996 40292
rect 15820 39564 15876 39620
rect 16268 39676 16324 39732
rect 15372 38556 15428 38612
rect 16604 39618 16660 39620
rect 16604 39566 16606 39618
rect 16606 39566 16658 39618
rect 16658 39566 16660 39618
rect 16604 39564 16660 39566
rect 16156 38162 16212 38164
rect 16156 38110 16158 38162
rect 16158 38110 16210 38162
rect 16210 38110 16212 38162
rect 16156 38108 16212 38110
rect 16940 39452 16996 39508
rect 17164 42364 17220 42420
rect 17388 43426 17444 43428
rect 17388 43374 17390 43426
rect 17390 43374 17442 43426
rect 17442 43374 17444 43426
rect 17388 43372 17444 43374
rect 17388 41970 17444 41972
rect 17388 41918 17390 41970
rect 17390 41918 17442 41970
rect 17442 41918 17444 41970
rect 17388 41916 17444 41918
rect 17724 44156 17780 44212
rect 17500 41804 17556 41860
rect 17612 43932 17668 43988
rect 17724 43708 17780 43764
rect 17388 41356 17444 41412
rect 17388 41186 17444 41188
rect 17388 41134 17390 41186
rect 17390 41134 17442 41186
rect 17442 41134 17444 41186
rect 17388 41132 17444 41134
rect 17276 41020 17332 41076
rect 17276 40684 17332 40740
rect 17388 40124 17444 40180
rect 17164 38780 17220 38836
rect 18172 46674 18228 46676
rect 18172 46622 18174 46674
rect 18174 46622 18226 46674
rect 18226 46622 18228 46674
rect 18172 46620 18228 46622
rect 18060 45388 18116 45444
rect 18284 45164 18340 45220
rect 18060 43932 18116 43988
rect 18732 50370 18788 50372
rect 18732 50318 18734 50370
rect 18734 50318 18786 50370
rect 18786 50318 18788 50370
rect 18732 50316 18788 50318
rect 18844 50092 18900 50148
rect 18732 49980 18788 50036
rect 19292 49810 19348 49812
rect 19292 49758 19294 49810
rect 19294 49758 19346 49810
rect 19346 49758 19348 49810
rect 19292 49756 19348 49758
rect 19180 49308 19236 49364
rect 18508 48748 18564 48804
rect 18732 48860 18788 48916
rect 19628 50594 19684 50596
rect 19628 50542 19630 50594
rect 19630 50542 19682 50594
rect 19682 50542 19684 50594
rect 19628 50540 19684 50542
rect 20300 52162 20356 52164
rect 20300 52110 20302 52162
rect 20302 52110 20354 52162
rect 20354 52110 20356 52162
rect 20300 52108 20356 52110
rect 20188 51324 20244 51380
rect 20412 51212 20468 51268
rect 20076 51154 20132 51156
rect 20076 51102 20078 51154
rect 20078 51102 20130 51154
rect 20130 51102 20132 51154
rect 20076 51100 20132 51102
rect 20748 52444 20804 52500
rect 20636 51938 20692 51940
rect 20636 51886 20638 51938
rect 20638 51886 20690 51938
rect 20690 51886 20692 51938
rect 20636 51884 20692 51886
rect 20860 51884 20916 51940
rect 20636 51436 20692 51492
rect 20748 51378 20804 51380
rect 20748 51326 20750 51378
rect 20750 51326 20802 51378
rect 20802 51326 20804 51378
rect 20748 51324 20804 51326
rect 20636 50876 20692 50932
rect 20748 50482 20804 50484
rect 20748 50430 20750 50482
rect 20750 50430 20802 50482
rect 20802 50430 20804 50482
rect 20748 50428 20804 50430
rect 19628 50316 19684 50372
rect 18732 48188 18788 48244
rect 18620 47516 18676 47572
rect 18732 47964 18788 48020
rect 18956 47516 19012 47572
rect 18732 46956 18788 47012
rect 18844 47068 18900 47124
rect 18508 46844 18564 46900
rect 18732 46396 18788 46452
rect 18732 46060 18788 46116
rect 18956 45890 19012 45892
rect 18956 45838 18958 45890
rect 18958 45838 19010 45890
rect 19010 45838 19012 45890
rect 18956 45836 19012 45838
rect 19404 47292 19460 47348
rect 19516 47628 19572 47684
rect 19404 46844 19460 46900
rect 19404 45724 19460 45780
rect 19180 45612 19236 45668
rect 19068 44828 19124 44884
rect 18844 44434 18900 44436
rect 18844 44382 18846 44434
rect 18846 44382 18898 44434
rect 18898 44382 18900 44434
rect 18844 44380 18900 44382
rect 18396 43484 18452 43540
rect 18060 42812 18116 42868
rect 17836 41580 17892 41636
rect 17948 41356 18004 41412
rect 18956 43820 19012 43876
rect 19964 50370 20020 50372
rect 19964 50318 19966 50370
rect 19966 50318 20018 50370
rect 20018 50318 20020 50370
rect 19964 50316 20020 50318
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 20524 50204 20580 50260
rect 20188 49922 20244 49924
rect 20188 49870 20190 49922
rect 20190 49870 20242 49922
rect 20242 49870 20244 49922
rect 20188 49868 20244 49870
rect 20412 49756 20468 49812
rect 19964 49698 20020 49700
rect 19964 49646 19966 49698
rect 19966 49646 20018 49698
rect 20018 49646 20020 49698
rect 19964 49644 20020 49646
rect 19852 49420 19908 49476
rect 20188 49138 20244 49140
rect 20188 49086 20190 49138
rect 20190 49086 20242 49138
rect 20242 49086 20244 49138
rect 20188 49084 20244 49086
rect 19964 49026 20020 49028
rect 19964 48974 19966 49026
rect 19966 48974 20018 49026
rect 20018 48974 20020 49026
rect 19964 48972 20020 48974
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 20300 48636 20356 48692
rect 20076 48242 20132 48244
rect 20076 48190 20078 48242
rect 20078 48190 20130 48242
rect 20130 48190 20132 48242
rect 20076 48188 20132 48190
rect 20188 48076 20244 48132
rect 19852 47628 19908 47684
rect 20300 47628 20356 47684
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 20412 47180 20468 47236
rect 20188 46396 20244 46452
rect 20300 46172 20356 46228
rect 19740 46060 19796 46116
rect 20412 46060 20468 46116
rect 19740 45778 19796 45780
rect 19740 45726 19742 45778
rect 19742 45726 19794 45778
rect 19794 45726 19796 45778
rect 19740 45724 19796 45726
rect 20636 48972 20692 49028
rect 20636 48018 20692 48020
rect 20636 47966 20638 48018
rect 20638 47966 20690 48018
rect 20690 47966 20692 48018
rect 20636 47964 20692 47966
rect 20748 47570 20804 47572
rect 20748 47518 20750 47570
rect 20750 47518 20802 47570
rect 20802 47518 20804 47570
rect 20748 47516 20804 47518
rect 20748 47180 20804 47236
rect 20076 45612 20132 45668
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 19628 45276 19684 45332
rect 19740 45164 19796 45220
rect 19292 44716 19348 44772
rect 18732 42978 18788 42980
rect 18732 42926 18734 42978
rect 18734 42926 18786 42978
rect 18786 42926 18788 42978
rect 18732 42924 18788 42926
rect 18284 42866 18340 42868
rect 18284 42814 18286 42866
rect 18286 42814 18338 42866
rect 18338 42814 18340 42866
rect 18284 42812 18340 42814
rect 18732 42754 18788 42756
rect 18732 42702 18734 42754
rect 18734 42702 18786 42754
rect 18786 42702 18788 42754
rect 18732 42700 18788 42702
rect 18956 42028 19012 42084
rect 18284 41244 18340 41300
rect 18396 41804 18452 41860
rect 17164 38108 17220 38164
rect 17724 41020 17780 41076
rect 17724 40460 17780 40516
rect 16268 37996 16324 38052
rect 15484 37772 15540 37828
rect 14028 37378 14084 37380
rect 14028 37326 14030 37378
rect 14030 37326 14082 37378
rect 14082 37326 14084 37378
rect 14028 37324 14084 37326
rect 15148 37378 15204 37380
rect 15148 37326 15150 37378
rect 15150 37326 15202 37378
rect 15202 37326 15204 37378
rect 15148 37324 15204 37326
rect 13132 36652 13188 36708
rect 13468 36540 13524 36596
rect 13580 36428 13636 36484
rect 12908 36204 12964 36260
rect 11116 35698 11172 35700
rect 11116 35646 11118 35698
rect 11118 35646 11170 35698
rect 11170 35646 11172 35698
rect 11116 35644 11172 35646
rect 13580 35810 13636 35812
rect 13580 35758 13582 35810
rect 13582 35758 13634 35810
rect 13634 35758 13636 35810
rect 13580 35756 13636 35758
rect 14588 36876 14644 36932
rect 11900 35644 11956 35700
rect 13244 35698 13300 35700
rect 13244 35646 13246 35698
rect 13246 35646 13298 35698
rect 13298 35646 13300 35698
rect 13244 35644 13300 35646
rect 13692 35644 13748 35700
rect 13916 36706 13972 36708
rect 13916 36654 13918 36706
rect 13918 36654 13970 36706
rect 13970 36654 13972 36706
rect 13916 36652 13972 36654
rect 12460 35586 12516 35588
rect 12460 35534 12462 35586
rect 12462 35534 12514 35586
rect 12514 35534 12516 35586
rect 12460 35532 12516 35534
rect 12012 35308 12068 35364
rect 12908 35026 12964 35028
rect 12908 34974 12910 35026
rect 12910 34974 12962 35026
rect 12962 34974 12964 35026
rect 12908 34972 12964 34974
rect 13468 34972 13524 35028
rect 11116 34748 11172 34804
rect 9996 34300 10052 34356
rect 8988 34076 9044 34132
rect 9548 33964 9604 34020
rect 5964 30098 6020 30100
rect 5964 30046 5966 30098
rect 5966 30046 6018 30098
rect 6018 30046 6020 30098
rect 5964 30044 6020 30046
rect 7868 30044 7924 30100
rect 7196 29820 7252 29876
rect 5068 29036 5124 29092
rect 5964 28700 6020 28756
rect 1932 27580 1988 27636
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 1708 26908 1764 26964
rect 4844 26908 4900 26964
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 2156 25564 2212 25620
rect 1708 24498 1764 24500
rect 1708 24446 1710 24498
rect 1710 24446 1762 24498
rect 1762 24446 1764 24498
rect 1708 24444 1764 24446
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 6972 28642 7028 28644
rect 6972 28590 6974 28642
rect 6974 28590 7026 28642
rect 7026 28590 7028 28642
rect 6972 28588 7028 28590
rect 6636 28476 6692 28532
rect 6076 27020 6132 27076
rect 7756 28700 7812 28756
rect 7644 28588 7700 28644
rect 7308 27580 7364 27636
rect 7308 27074 7364 27076
rect 7308 27022 7310 27074
rect 7310 27022 7362 27074
rect 7362 27022 7364 27074
rect 7308 27020 7364 27022
rect 8764 30156 8820 30212
rect 8540 30098 8596 30100
rect 8540 30046 8542 30098
rect 8542 30046 8594 30098
rect 8594 30046 8596 30098
rect 8540 30044 8596 30046
rect 8428 28476 8484 28532
rect 10556 34412 10612 34468
rect 15372 36876 15428 36932
rect 14924 36652 14980 36708
rect 14140 36092 14196 36148
rect 14252 35922 14308 35924
rect 14252 35870 14254 35922
rect 14254 35870 14306 35922
rect 14306 35870 14308 35922
rect 14252 35868 14308 35870
rect 14140 35698 14196 35700
rect 14140 35646 14142 35698
rect 14142 35646 14194 35698
rect 14194 35646 14196 35698
rect 14140 35644 14196 35646
rect 14812 35698 14868 35700
rect 14812 35646 14814 35698
rect 14814 35646 14866 35698
rect 14866 35646 14868 35698
rect 14812 35644 14868 35646
rect 14028 35196 14084 35252
rect 11340 34690 11396 34692
rect 11340 34638 11342 34690
rect 11342 34638 11394 34690
rect 11394 34638 11396 34690
rect 11340 34636 11396 34638
rect 11116 33628 11172 33684
rect 13020 33628 13076 33684
rect 11676 33346 11732 33348
rect 11676 33294 11678 33346
rect 11678 33294 11730 33346
rect 11730 33294 11732 33346
rect 11676 33292 11732 33294
rect 10892 32732 10948 32788
rect 12012 33068 12068 33124
rect 10108 31724 10164 31780
rect 12572 33122 12628 33124
rect 12572 33070 12574 33122
rect 12574 33070 12626 33122
rect 12626 33070 12628 33122
rect 12572 33068 12628 33070
rect 9100 29820 9156 29876
rect 9884 30044 9940 30100
rect 11228 30210 11284 30212
rect 11228 30158 11230 30210
rect 11230 30158 11282 30210
rect 11282 30158 11284 30210
rect 11228 30156 11284 30158
rect 14476 34972 14532 35028
rect 14252 34412 14308 34468
rect 15932 37490 15988 37492
rect 15932 37438 15934 37490
rect 15934 37438 15986 37490
rect 15986 37438 15988 37490
rect 15932 37436 15988 37438
rect 15596 37266 15652 37268
rect 15596 37214 15598 37266
rect 15598 37214 15650 37266
rect 15650 37214 15652 37266
rect 15596 37212 15652 37214
rect 16604 36876 16660 36932
rect 15372 35756 15428 35812
rect 16268 35922 16324 35924
rect 16268 35870 16270 35922
rect 16270 35870 16322 35922
rect 16322 35870 16324 35922
rect 16268 35868 16324 35870
rect 15372 34860 15428 34916
rect 17052 36092 17108 36148
rect 17388 36092 17444 36148
rect 17500 38444 17556 38500
rect 17612 37490 17668 37492
rect 17612 37438 17614 37490
rect 17614 37438 17666 37490
rect 17666 37438 17668 37490
rect 17612 37436 17668 37438
rect 17836 40236 17892 40292
rect 17836 39452 17892 39508
rect 17948 39564 18004 39620
rect 17948 38834 18004 38836
rect 17948 38782 17950 38834
rect 17950 38782 18002 38834
rect 18002 38782 18004 38834
rect 17948 38780 18004 38782
rect 17836 38050 17892 38052
rect 17836 37998 17838 38050
rect 17838 37998 17890 38050
rect 17890 37998 17892 38050
rect 17836 37996 17892 37998
rect 17948 37772 18004 37828
rect 18396 41132 18452 41188
rect 18956 41244 19012 41300
rect 20188 45218 20244 45220
rect 20188 45166 20190 45218
rect 20190 45166 20242 45218
rect 20242 45166 20244 45218
rect 20188 45164 20244 45166
rect 19964 45052 20020 45108
rect 19404 43596 19460 43652
rect 19516 44492 19572 44548
rect 19516 44268 19572 44324
rect 19852 44322 19908 44324
rect 19852 44270 19854 44322
rect 19854 44270 19906 44322
rect 19906 44270 19908 44322
rect 19852 44268 19908 44270
rect 19964 44210 20020 44212
rect 19964 44158 19966 44210
rect 19966 44158 20018 44210
rect 20018 44158 20020 44210
rect 19964 44156 20020 44158
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 19740 43596 19796 43652
rect 19740 43372 19796 43428
rect 18844 40796 18900 40852
rect 19404 42642 19460 42644
rect 19404 42590 19406 42642
rect 19406 42590 19458 42642
rect 19458 42590 19460 42642
rect 19404 42588 19460 42590
rect 21868 56194 21924 56196
rect 21868 56142 21870 56194
rect 21870 56142 21922 56194
rect 21922 56142 21924 56194
rect 21868 56140 21924 56142
rect 22652 56140 22708 56196
rect 21308 56082 21364 56084
rect 21308 56030 21310 56082
rect 21310 56030 21362 56082
rect 21362 56030 21364 56082
rect 21308 56028 21364 56030
rect 21756 55804 21812 55860
rect 22540 55580 22596 55636
rect 22428 55356 22484 55412
rect 22204 55186 22260 55188
rect 22204 55134 22206 55186
rect 22206 55134 22258 55186
rect 22258 55134 22260 55186
rect 22204 55132 22260 55134
rect 21756 54572 21812 54628
rect 22764 55580 22820 55636
rect 22652 54738 22708 54740
rect 22652 54686 22654 54738
rect 22654 54686 22706 54738
rect 22706 54686 22708 54738
rect 22652 54684 22708 54686
rect 21196 53900 21252 53956
rect 22092 54236 22148 54292
rect 21308 52946 21364 52948
rect 21308 52894 21310 52946
rect 21310 52894 21362 52946
rect 21362 52894 21364 52946
rect 21308 52892 21364 52894
rect 21644 52780 21700 52836
rect 21420 52444 21476 52500
rect 21420 52220 21476 52276
rect 21084 52108 21140 52164
rect 21644 52108 21700 52164
rect 21196 51772 21252 51828
rect 21196 51378 21252 51380
rect 21196 51326 21198 51378
rect 21198 51326 21250 51378
rect 21250 51326 21252 51378
rect 21196 51324 21252 51326
rect 21868 51602 21924 51604
rect 21868 51550 21870 51602
rect 21870 51550 21922 51602
rect 21922 51550 21924 51602
rect 21868 51548 21924 51550
rect 21756 51436 21812 51492
rect 21084 50428 21140 50484
rect 21196 50652 21252 50708
rect 20972 48972 21028 49028
rect 21084 49868 21140 49924
rect 20972 47068 21028 47124
rect 21420 50316 21476 50372
rect 21308 49532 21364 49588
rect 21308 48972 21364 49028
rect 21644 51212 21700 51268
rect 21644 50316 21700 50372
rect 21644 49532 21700 49588
rect 21644 47628 21700 47684
rect 21756 48188 21812 48244
rect 21084 46732 21140 46788
rect 20860 45948 20916 46004
rect 20524 44828 20580 44884
rect 20524 44210 20580 44212
rect 20524 44158 20526 44210
rect 20526 44158 20578 44210
rect 20578 44158 20580 44210
rect 20524 44156 20580 44158
rect 20412 43596 20468 43652
rect 20412 42924 20468 42980
rect 20748 44044 20804 44100
rect 20972 45500 21028 45556
rect 21308 46060 21364 46116
rect 21196 44994 21252 44996
rect 21196 44942 21198 44994
rect 21198 44942 21250 44994
rect 21250 44942 21252 44994
rect 21196 44940 21252 44942
rect 21308 44322 21364 44324
rect 21308 44270 21310 44322
rect 21310 44270 21362 44322
rect 21362 44270 21364 44322
rect 21308 44268 21364 44270
rect 21084 43650 21140 43652
rect 21084 43598 21086 43650
rect 21086 43598 21138 43650
rect 21138 43598 21140 43650
rect 21084 43596 21140 43598
rect 20860 43260 20916 43316
rect 19292 42028 19348 42084
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 20860 42812 20916 42868
rect 19964 42082 20020 42084
rect 19964 42030 19966 42082
rect 19966 42030 20018 42082
rect 20018 42030 20020 42082
rect 19964 42028 20020 42030
rect 19404 41970 19460 41972
rect 19404 41918 19406 41970
rect 19406 41918 19458 41970
rect 19458 41918 19460 41970
rect 19404 41916 19460 41918
rect 19740 41970 19796 41972
rect 19740 41918 19742 41970
rect 19742 41918 19794 41970
rect 19794 41918 19796 41970
rect 19740 41916 19796 41918
rect 19292 41356 19348 41412
rect 19292 41020 19348 41076
rect 18956 40236 19012 40292
rect 18956 39900 19012 39956
rect 18396 39676 18452 39732
rect 18284 39340 18340 39396
rect 18956 39340 19012 39396
rect 18508 37884 18564 37940
rect 17500 35756 17556 35812
rect 18284 36764 18340 36820
rect 17724 36258 17780 36260
rect 17724 36206 17726 36258
rect 17726 36206 17778 36258
rect 17778 36206 17780 36258
rect 17724 36204 17780 36206
rect 16380 34748 16436 34804
rect 16828 35196 16884 35252
rect 14700 34412 14756 34468
rect 18396 36370 18452 36372
rect 18396 36318 18398 36370
rect 18398 36318 18450 36370
rect 18450 36318 18452 36370
rect 18396 36316 18452 36318
rect 17836 34972 17892 35028
rect 18396 34802 18452 34804
rect 18396 34750 18398 34802
rect 18398 34750 18450 34802
rect 18450 34750 18452 34802
rect 18396 34748 18452 34750
rect 18732 37490 18788 37492
rect 18732 37438 18734 37490
rect 18734 37438 18786 37490
rect 18786 37438 18788 37490
rect 18732 37436 18788 37438
rect 19180 40348 19236 40404
rect 19292 39618 19348 39620
rect 19292 39566 19294 39618
rect 19294 39566 19346 39618
rect 19346 39566 19348 39618
rect 19292 39564 19348 39566
rect 19180 39228 19236 39284
rect 19628 41356 19684 41412
rect 20188 41580 20244 41636
rect 19628 41074 19684 41076
rect 19628 41022 19630 41074
rect 19630 41022 19682 41074
rect 19682 41022 19684 41074
rect 19628 41020 19684 41022
rect 20076 40962 20132 40964
rect 20076 40910 20078 40962
rect 20078 40910 20130 40962
rect 20130 40910 20132 40962
rect 20076 40908 20132 40910
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 19740 40572 19796 40628
rect 19740 39506 19796 39508
rect 19740 39454 19742 39506
rect 19742 39454 19794 39506
rect 19794 39454 19796 39506
rect 19740 39452 19796 39454
rect 19516 39228 19572 39284
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19068 38556 19124 38612
rect 19964 38722 20020 38724
rect 19964 38670 19966 38722
rect 19966 38670 20018 38722
rect 20018 38670 20020 38722
rect 19964 38668 20020 38670
rect 19292 38162 19348 38164
rect 19292 38110 19294 38162
rect 19294 38110 19346 38162
rect 19346 38110 19348 38162
rect 19292 38108 19348 38110
rect 19628 37996 19684 38052
rect 18844 36764 18900 36820
rect 18956 36428 19012 36484
rect 20524 41020 20580 41076
rect 20188 37826 20244 37828
rect 20188 37774 20190 37826
rect 20190 37774 20242 37826
rect 20242 37774 20244 37826
rect 20188 37772 20244 37774
rect 20300 38556 20356 38612
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19404 36428 19460 36484
rect 19852 37100 19908 37156
rect 20188 37212 20244 37268
rect 20748 41020 20804 41076
rect 20748 40796 20804 40852
rect 20748 40626 20804 40628
rect 20748 40574 20750 40626
rect 20750 40574 20802 40626
rect 20802 40574 20804 40626
rect 20748 40572 20804 40574
rect 20636 39788 20692 39844
rect 20748 40012 20804 40068
rect 20748 39228 20804 39284
rect 20860 38946 20916 38948
rect 20860 38894 20862 38946
rect 20862 38894 20914 38946
rect 20914 38894 20916 38946
rect 20860 38892 20916 38894
rect 20636 38610 20692 38612
rect 20636 38558 20638 38610
rect 20638 38558 20690 38610
rect 20690 38558 20692 38610
rect 20636 38556 20692 38558
rect 20748 38050 20804 38052
rect 20748 37998 20750 38050
rect 20750 37998 20802 38050
rect 20802 37998 20804 38050
rect 20748 37996 20804 37998
rect 20524 37100 20580 37156
rect 20188 36540 20244 36596
rect 19516 36092 19572 36148
rect 18620 34860 18676 34916
rect 14140 33964 14196 34020
rect 13692 33180 13748 33236
rect 13580 33122 13636 33124
rect 13580 33070 13582 33122
rect 13582 33070 13634 33122
rect 13634 33070 13636 33122
rect 13580 33068 13636 33070
rect 15260 34018 15316 34020
rect 15260 33966 15262 34018
rect 15262 33966 15314 34018
rect 15314 33966 15316 34018
rect 15260 33964 15316 33966
rect 14028 33068 14084 33124
rect 14588 33516 14644 33572
rect 18396 33964 18452 34020
rect 18508 33740 18564 33796
rect 19068 34412 19124 34468
rect 17164 33404 17220 33460
rect 15260 33292 15316 33348
rect 16604 33292 16660 33348
rect 18732 33516 18788 33572
rect 19292 35196 19348 35252
rect 17500 33346 17556 33348
rect 17500 33294 17502 33346
rect 17502 33294 17554 33346
rect 17554 33294 17556 33346
rect 17500 33292 17556 33294
rect 19404 34914 19460 34916
rect 19404 34862 19406 34914
rect 19406 34862 19458 34914
rect 19458 34862 19460 34914
rect 19404 34860 19460 34862
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19852 35922 19908 35924
rect 19852 35870 19854 35922
rect 19854 35870 19906 35922
rect 19906 35870 19908 35922
rect 19852 35868 19908 35870
rect 20412 35698 20468 35700
rect 20412 35646 20414 35698
rect 20414 35646 20466 35698
rect 20466 35646 20468 35698
rect 20412 35644 20468 35646
rect 20076 35196 20132 35252
rect 19628 34972 19684 35028
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19516 34300 19572 34356
rect 19852 34300 19908 34356
rect 19628 34242 19684 34244
rect 19628 34190 19630 34242
rect 19630 34190 19682 34242
rect 19682 34190 19684 34242
rect 19628 34188 19684 34190
rect 19516 34130 19572 34132
rect 19516 34078 19518 34130
rect 19518 34078 19570 34130
rect 19570 34078 19572 34130
rect 19516 34076 19572 34078
rect 18956 33122 19012 33124
rect 18956 33070 18958 33122
rect 18958 33070 19010 33122
rect 19010 33070 19012 33122
rect 18956 33068 19012 33070
rect 18508 32620 18564 32676
rect 11788 30210 11844 30212
rect 11788 30158 11790 30210
rect 11790 30158 11842 30210
rect 11842 30158 11844 30210
rect 11788 30156 11844 30158
rect 10780 30044 10836 30100
rect 9772 29314 9828 29316
rect 9772 29262 9774 29314
rect 9774 29262 9826 29314
rect 9826 29262 9828 29314
rect 9772 29260 9828 29262
rect 11004 29426 11060 29428
rect 11004 29374 11006 29426
rect 11006 29374 11058 29426
rect 11058 29374 11060 29426
rect 11004 29372 11060 29374
rect 10444 29260 10500 29316
rect 9212 28588 9268 28644
rect 9100 28364 9156 28420
rect 8428 27970 8484 27972
rect 8428 27918 8430 27970
rect 8430 27918 8482 27970
rect 8482 27918 8484 27970
rect 8428 27916 8484 27918
rect 8092 27634 8148 27636
rect 8092 27582 8094 27634
rect 8094 27582 8146 27634
rect 8146 27582 8148 27634
rect 8092 27580 8148 27582
rect 7532 27020 7588 27076
rect 6860 26178 6916 26180
rect 6860 26126 6862 26178
rect 6862 26126 6914 26178
rect 6914 26126 6916 26178
rect 6860 26124 6916 26126
rect 6412 25788 6468 25844
rect 5964 25506 6020 25508
rect 5964 25454 5966 25506
rect 5966 25454 6018 25506
rect 6018 25454 6020 25506
rect 5964 25452 6020 25454
rect 5628 25394 5684 25396
rect 5628 25342 5630 25394
rect 5630 25342 5682 25394
rect 5682 25342 5684 25394
rect 5628 25340 5684 25342
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 1708 20860 1764 20916
rect 5628 22876 5684 22932
rect 7420 26012 7476 26068
rect 6860 25394 6916 25396
rect 6860 25342 6862 25394
rect 6862 25342 6914 25394
rect 6914 25342 6916 25394
rect 6860 25340 6916 25342
rect 6636 24610 6692 24612
rect 6636 24558 6638 24610
rect 6638 24558 6690 24610
rect 6690 24558 6692 24610
rect 6636 24556 6692 24558
rect 6076 22370 6132 22372
rect 6076 22318 6078 22370
rect 6078 22318 6130 22370
rect 6130 22318 6132 22370
rect 6076 22316 6132 22318
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4396 17836 4452 17892
rect 1708 17554 1764 17556
rect 1708 17502 1710 17554
rect 1710 17502 1762 17554
rect 1762 17502 1764 17554
rect 1708 17500 1764 17502
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 5852 20018 5908 20020
rect 5852 19966 5854 20018
rect 5854 19966 5906 20018
rect 5906 19966 5908 20018
rect 5852 19964 5908 19966
rect 5964 18620 6020 18676
rect 6076 18450 6132 18452
rect 6076 18398 6078 18450
rect 6078 18398 6130 18450
rect 6130 18398 6132 18450
rect 6076 18396 6132 18398
rect 5068 17666 5124 17668
rect 5068 17614 5070 17666
rect 5070 17614 5122 17666
rect 5122 17614 5124 17666
rect 5068 17612 5124 17614
rect 5740 17666 5796 17668
rect 5740 17614 5742 17666
rect 5742 17614 5794 17666
rect 5794 17614 5796 17666
rect 5740 17612 5796 17614
rect 6076 17164 6132 17220
rect 5516 17106 5572 17108
rect 5516 17054 5518 17106
rect 5518 17054 5570 17106
rect 5570 17054 5572 17106
rect 5516 17052 5572 17054
rect 7308 23938 7364 23940
rect 7308 23886 7310 23938
rect 7310 23886 7362 23938
rect 7362 23886 7364 23938
rect 7308 23884 7364 23886
rect 7196 22876 7252 22932
rect 6524 21868 6580 21924
rect 6524 21644 6580 21700
rect 6300 20690 6356 20692
rect 6300 20638 6302 20690
rect 6302 20638 6354 20690
rect 6354 20638 6356 20690
rect 6300 20636 6356 20638
rect 6972 22370 7028 22372
rect 6972 22318 6974 22370
rect 6974 22318 7026 22370
rect 7026 22318 7028 22370
rect 6972 22316 7028 22318
rect 6636 21532 6692 21588
rect 6748 22092 6804 22148
rect 8092 25452 8148 25508
rect 8540 27244 8596 27300
rect 7868 24668 7924 24724
rect 8652 25452 8708 25508
rect 8540 24722 8596 24724
rect 8540 24670 8542 24722
rect 8542 24670 8594 24722
rect 8594 24670 8596 24722
rect 8540 24668 8596 24670
rect 8204 23884 8260 23940
rect 7420 22316 7476 22372
rect 7532 22092 7588 22148
rect 6972 20188 7028 20244
rect 6524 18508 6580 18564
rect 7084 20018 7140 20020
rect 7084 19966 7086 20018
rect 7086 19966 7138 20018
rect 7138 19966 7140 20018
rect 7084 19964 7140 19966
rect 7084 19292 7140 19348
rect 6748 19180 6804 19236
rect 6748 18396 6804 18452
rect 4956 16380 5012 16436
rect 4732 15986 4788 15988
rect 4732 15934 4734 15986
rect 4734 15934 4786 15986
rect 4786 15934 4788 15986
rect 4732 15932 4788 15934
rect 5068 15538 5124 15540
rect 5068 15486 5070 15538
rect 5070 15486 5122 15538
rect 5122 15486 5124 15538
rect 5068 15484 5124 15486
rect 5516 16380 5572 16436
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 5180 14642 5236 14644
rect 5180 14590 5182 14642
rect 5182 14590 5234 14642
rect 5234 14590 5236 14642
rect 5180 14588 5236 14590
rect 5964 15596 6020 15652
rect 5852 14812 5908 14868
rect 6860 17948 6916 18004
rect 7084 19122 7140 19124
rect 7084 19070 7086 19122
rect 7086 19070 7138 19122
rect 7138 19070 7140 19122
rect 7084 19068 7140 19070
rect 6972 17276 7028 17332
rect 7308 21586 7364 21588
rect 7308 21534 7310 21586
rect 7310 21534 7362 21586
rect 7362 21534 7364 21586
rect 7308 21532 7364 21534
rect 7308 20076 7364 20132
rect 7532 19964 7588 20020
rect 7308 19180 7364 19236
rect 8092 21532 8148 21588
rect 7868 21420 7924 21476
rect 7980 20188 8036 20244
rect 7756 19292 7812 19348
rect 8092 19964 8148 20020
rect 7308 17612 7364 17668
rect 7084 17052 7140 17108
rect 6860 16940 6916 16996
rect 7420 17052 7476 17108
rect 6748 16828 6804 16884
rect 6636 16268 6692 16324
rect 5852 14588 5908 14644
rect 6636 14924 6692 14980
rect 5404 14364 5460 14420
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 6188 14530 6244 14532
rect 6188 14478 6190 14530
rect 6190 14478 6242 14530
rect 6242 14478 6244 14530
rect 6188 14476 6244 14478
rect 6524 14364 6580 14420
rect 6188 13020 6244 13076
rect 6636 13746 6692 13748
rect 6636 13694 6638 13746
rect 6638 13694 6690 13746
rect 6690 13694 6692 13746
rect 6636 13692 6692 13694
rect 6748 12796 6804 12852
rect 7420 16380 7476 16436
rect 7532 16098 7588 16100
rect 7532 16046 7534 16098
rect 7534 16046 7586 16098
rect 7586 16046 7588 16098
rect 7532 16044 7588 16046
rect 8540 22370 8596 22372
rect 8540 22318 8542 22370
rect 8542 22318 8594 22370
rect 8594 22318 8596 22370
rect 8540 22316 8596 22318
rect 8428 21644 8484 21700
rect 9548 27970 9604 27972
rect 9548 27918 9550 27970
rect 9550 27918 9602 27970
rect 9602 27918 9604 27970
rect 9548 27916 9604 27918
rect 10108 28642 10164 28644
rect 10108 28590 10110 28642
rect 10110 28590 10162 28642
rect 10162 28590 10164 28642
rect 10108 28588 10164 28590
rect 9884 27970 9940 27972
rect 9884 27918 9886 27970
rect 9886 27918 9938 27970
rect 9938 27918 9940 27970
rect 9884 27916 9940 27918
rect 9772 27804 9828 27860
rect 11004 29148 11060 29204
rect 10556 28700 10612 28756
rect 10892 27916 10948 27972
rect 10444 27356 10500 27412
rect 8988 26962 9044 26964
rect 8988 26910 8990 26962
rect 8990 26910 9042 26962
rect 9042 26910 9044 26962
rect 8988 26908 9044 26910
rect 9548 27186 9604 27188
rect 9548 27134 9550 27186
rect 9550 27134 9602 27186
rect 9602 27134 9604 27186
rect 9548 27132 9604 27134
rect 9436 26236 9492 26292
rect 9324 25730 9380 25732
rect 9324 25678 9326 25730
rect 9326 25678 9378 25730
rect 9378 25678 9380 25730
rect 9324 25676 9380 25678
rect 9324 25452 9380 25508
rect 8988 25116 9044 25172
rect 10444 27074 10500 27076
rect 10444 27022 10446 27074
rect 10446 27022 10498 27074
rect 10498 27022 10500 27074
rect 10444 27020 10500 27022
rect 10780 27858 10836 27860
rect 10780 27806 10782 27858
rect 10782 27806 10834 27858
rect 10834 27806 10836 27858
rect 10780 27804 10836 27806
rect 10108 26290 10164 26292
rect 10108 26238 10110 26290
rect 10110 26238 10162 26290
rect 10162 26238 10164 26290
rect 10108 26236 10164 26238
rect 13916 30380 13972 30436
rect 13692 30210 13748 30212
rect 13692 30158 13694 30210
rect 13694 30158 13746 30210
rect 13746 30158 13748 30210
rect 13692 30156 13748 30158
rect 17500 31500 17556 31556
rect 18172 31554 18228 31556
rect 18172 31502 18174 31554
rect 18174 31502 18226 31554
rect 18226 31502 18228 31554
rect 18172 31500 18228 31502
rect 17836 31164 17892 31220
rect 16716 31052 16772 31108
rect 15484 30380 15540 30436
rect 17052 30492 17108 30548
rect 16940 30098 16996 30100
rect 16940 30046 16942 30098
rect 16942 30046 16994 30098
rect 16994 30046 16996 30098
rect 16940 30044 16996 30046
rect 12460 29148 12516 29204
rect 12012 28812 12068 28868
rect 13468 28812 13524 28868
rect 13916 28642 13972 28644
rect 13916 28590 13918 28642
rect 13918 28590 13970 28642
rect 13970 28590 13972 28642
rect 13916 28588 13972 28590
rect 11228 27916 11284 27972
rect 11228 27468 11284 27524
rect 10892 27020 10948 27076
rect 11004 27356 11060 27412
rect 10668 26236 10724 26292
rect 11116 27244 11172 27300
rect 10556 25676 10612 25732
rect 9884 25506 9940 25508
rect 9884 25454 9886 25506
rect 9886 25454 9938 25506
rect 9938 25454 9940 25506
rect 9884 25452 9940 25454
rect 9884 25228 9940 25284
rect 8988 24834 9044 24836
rect 8988 24782 8990 24834
rect 8990 24782 9042 24834
rect 9042 24782 9044 24834
rect 8988 24780 9044 24782
rect 9548 24722 9604 24724
rect 9548 24670 9550 24722
rect 9550 24670 9602 24722
rect 9602 24670 9604 24722
rect 9548 24668 9604 24670
rect 9324 23100 9380 23156
rect 9996 23826 10052 23828
rect 9996 23774 9998 23826
rect 9998 23774 10050 23826
rect 10050 23774 10052 23826
rect 9996 23772 10052 23774
rect 9884 22428 9940 22484
rect 8988 22370 9044 22372
rect 8988 22318 8990 22370
rect 8990 22318 9042 22370
rect 9042 22318 9044 22370
rect 8988 22316 9044 22318
rect 8988 21474 9044 21476
rect 8988 21422 8990 21474
rect 8990 21422 9042 21474
rect 9042 21422 9044 21474
rect 8988 21420 9044 21422
rect 8316 20748 8372 20804
rect 8652 20524 8708 20580
rect 8540 20018 8596 20020
rect 8540 19966 8542 20018
rect 8542 19966 8594 20018
rect 8594 19966 8596 20018
rect 8540 19964 8596 19966
rect 7980 18620 8036 18676
rect 8316 18562 8372 18564
rect 8316 18510 8318 18562
rect 8318 18510 8370 18562
rect 8370 18510 8372 18562
rect 8316 18508 8372 18510
rect 7756 17778 7812 17780
rect 7756 17726 7758 17778
rect 7758 17726 7810 17778
rect 7810 17726 7812 17778
rect 7756 17724 7812 17726
rect 7756 17106 7812 17108
rect 7756 17054 7758 17106
rect 7758 17054 7810 17106
rect 7810 17054 7812 17106
rect 7756 17052 7812 17054
rect 7756 16828 7812 16884
rect 7308 15260 7364 15316
rect 7196 14588 7252 14644
rect 7420 14252 7476 14308
rect 7644 15148 7700 15204
rect 8092 17724 8148 17780
rect 8764 19794 8820 19796
rect 8764 19742 8766 19794
rect 8766 19742 8818 19794
rect 8818 19742 8820 19794
rect 8764 19740 8820 19742
rect 9324 20748 9380 20804
rect 9772 21084 9828 21140
rect 9212 20412 9268 20468
rect 9100 19234 9156 19236
rect 9100 19182 9102 19234
rect 9102 19182 9154 19234
rect 9154 19182 9156 19234
rect 9100 19180 9156 19182
rect 8652 18956 8708 19012
rect 8988 18844 9044 18900
rect 8988 18620 9044 18676
rect 8876 18508 8932 18564
rect 8428 17724 8484 17780
rect 8652 17836 8708 17892
rect 8316 17666 8372 17668
rect 8316 17614 8318 17666
rect 8318 17614 8370 17666
rect 8370 17614 8372 17666
rect 8316 17612 8372 17614
rect 8092 15708 8148 15764
rect 8652 16994 8708 16996
rect 8652 16942 8654 16994
rect 8654 16942 8706 16994
rect 8706 16942 8708 16994
rect 8652 16940 8708 16942
rect 8876 16156 8932 16212
rect 7868 14588 7924 14644
rect 7756 13970 7812 13972
rect 7756 13918 7758 13970
rect 7758 13918 7810 13970
rect 7810 13918 7812 13970
rect 7756 13916 7812 13918
rect 6972 12962 7028 12964
rect 6972 12910 6974 12962
rect 6974 12910 7026 12962
rect 7026 12910 7028 12962
rect 6972 12908 7028 12910
rect 7308 12850 7364 12852
rect 7308 12798 7310 12850
rect 7310 12798 7362 12850
rect 7362 12798 7364 12850
rect 7308 12796 7364 12798
rect 7308 12348 7364 12404
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 6636 11564 6692 11620
rect 7084 11452 7140 11508
rect 7868 13356 7924 13412
rect 8764 15372 8820 15428
rect 8316 14642 8372 14644
rect 8316 14590 8318 14642
rect 8318 14590 8370 14642
rect 8370 14590 8372 14642
rect 8316 14588 8372 14590
rect 8316 13916 8372 13972
rect 8204 13580 8260 13636
rect 8652 14418 8708 14420
rect 8652 14366 8654 14418
rect 8654 14366 8706 14418
rect 8706 14366 8708 14418
rect 8652 14364 8708 14366
rect 9660 19234 9716 19236
rect 9660 19182 9662 19234
rect 9662 19182 9714 19234
rect 9714 19182 9716 19234
rect 9660 19180 9716 19182
rect 9884 19068 9940 19124
rect 9548 19010 9604 19012
rect 9548 18958 9550 19010
rect 9550 18958 9602 19010
rect 9602 18958 9604 19010
rect 9548 18956 9604 18958
rect 9436 18620 9492 18676
rect 9772 18508 9828 18564
rect 8876 13970 8932 13972
rect 8876 13918 8878 13970
rect 8878 13918 8930 13970
rect 8930 13918 8932 13970
rect 8876 13916 8932 13918
rect 9212 15932 9268 15988
rect 7868 11954 7924 11956
rect 7868 11902 7870 11954
rect 7870 11902 7922 11954
rect 7922 11902 7924 11954
rect 7868 11900 7924 11902
rect 7532 11676 7588 11732
rect 7756 11564 7812 11620
rect 8204 12402 8260 12404
rect 8204 12350 8206 12402
rect 8206 12350 8258 12402
rect 8258 12350 8260 12402
rect 8204 12348 8260 12350
rect 9100 13970 9156 13972
rect 9100 13918 9102 13970
rect 9102 13918 9154 13970
rect 9154 13918 9156 13970
rect 9100 13916 9156 13918
rect 8092 11340 8148 11396
rect 8652 12796 8708 12852
rect 8316 11676 8372 11732
rect 7420 10780 7476 10836
rect 8204 10834 8260 10836
rect 8204 10782 8206 10834
rect 8206 10782 8258 10834
rect 8258 10782 8260 10834
rect 8204 10780 8260 10782
rect 8764 12178 8820 12180
rect 8764 12126 8766 12178
rect 8766 12126 8818 12178
rect 8818 12126 8820 12178
rect 8764 12124 8820 12126
rect 9772 18338 9828 18340
rect 9772 18286 9774 18338
rect 9774 18286 9826 18338
rect 9826 18286 9828 18338
rect 9772 18284 9828 18286
rect 9772 18060 9828 18116
rect 9772 17276 9828 17332
rect 9660 16268 9716 16324
rect 9548 16044 9604 16100
rect 9324 14252 9380 14308
rect 9660 12348 9716 12404
rect 10108 22876 10164 22932
rect 10220 20802 10276 20804
rect 10220 20750 10222 20802
rect 10222 20750 10274 20802
rect 10274 20750 10276 20802
rect 10220 20748 10276 20750
rect 10108 20636 10164 20692
rect 10108 18284 10164 18340
rect 10220 19292 10276 19348
rect 9996 17500 10052 17556
rect 10108 17612 10164 17668
rect 9884 16044 9940 16100
rect 9996 16828 10052 16884
rect 11004 25506 11060 25508
rect 11004 25454 11006 25506
rect 11006 25454 11058 25506
rect 11058 25454 11060 25506
rect 11004 25452 11060 25454
rect 11004 24444 11060 24500
rect 11004 23324 11060 23380
rect 11004 23154 11060 23156
rect 11004 23102 11006 23154
rect 11006 23102 11058 23154
rect 11058 23102 11060 23154
rect 11004 23100 11060 23102
rect 10892 21474 10948 21476
rect 10892 21422 10894 21474
rect 10894 21422 10946 21474
rect 10946 21422 10948 21474
rect 10892 21420 10948 21422
rect 10780 20748 10836 20804
rect 12348 27916 12404 27972
rect 11676 27634 11732 27636
rect 11676 27582 11678 27634
rect 11678 27582 11730 27634
rect 11730 27582 11732 27634
rect 11676 27580 11732 27582
rect 12236 27132 12292 27188
rect 11564 27074 11620 27076
rect 11564 27022 11566 27074
rect 11566 27022 11618 27074
rect 11618 27022 11620 27074
rect 11564 27020 11620 27022
rect 12124 26962 12180 26964
rect 12124 26910 12126 26962
rect 12126 26910 12178 26962
rect 12178 26910 12180 26962
rect 12124 26908 12180 26910
rect 11340 25340 11396 25396
rect 11452 25452 11508 25508
rect 11452 24780 11508 24836
rect 11340 23212 11396 23268
rect 11340 21980 11396 22036
rect 12908 27074 12964 27076
rect 12908 27022 12910 27074
rect 12910 27022 12962 27074
rect 12962 27022 12964 27074
rect 12908 27020 12964 27022
rect 12460 26684 12516 26740
rect 12124 25900 12180 25956
rect 11676 25564 11732 25620
rect 11900 25676 11956 25732
rect 11788 25340 11844 25396
rect 12012 25228 12068 25284
rect 11900 24892 11956 24948
rect 11900 24556 11956 24612
rect 11788 23772 11844 23828
rect 11564 22876 11620 22932
rect 11676 23324 11732 23380
rect 11452 22764 11508 22820
rect 11676 22316 11732 22372
rect 11564 21868 11620 21924
rect 11676 21980 11732 22036
rect 11228 21756 11284 21812
rect 10668 19404 10724 19460
rect 11564 21698 11620 21700
rect 11564 21646 11566 21698
rect 11566 21646 11618 21698
rect 11618 21646 11620 21698
rect 11564 21644 11620 21646
rect 10556 18620 10612 18676
rect 10332 18562 10388 18564
rect 10332 18510 10334 18562
rect 10334 18510 10386 18562
rect 10386 18510 10388 18562
rect 10332 18508 10388 18510
rect 10444 18450 10500 18452
rect 10444 18398 10446 18450
rect 10446 18398 10498 18450
rect 10498 18398 10500 18450
rect 10444 18396 10500 18398
rect 10444 18172 10500 18228
rect 10332 17948 10388 18004
rect 10332 16940 10388 16996
rect 11004 19404 11060 19460
rect 10668 17500 10724 17556
rect 10444 15932 10500 15988
rect 10892 19122 10948 19124
rect 10892 19070 10894 19122
rect 10894 19070 10946 19122
rect 10946 19070 10948 19122
rect 10892 19068 10948 19070
rect 10780 15372 10836 15428
rect 10220 13746 10276 13748
rect 10220 13694 10222 13746
rect 10222 13694 10274 13746
rect 10274 13694 10276 13746
rect 10220 13692 10276 13694
rect 10332 13634 10388 13636
rect 10332 13582 10334 13634
rect 10334 13582 10386 13634
rect 10386 13582 10388 13634
rect 10332 13580 10388 13582
rect 10220 13468 10276 13524
rect 10108 13074 10164 13076
rect 10108 13022 10110 13074
rect 10110 13022 10162 13074
rect 10162 13022 10164 13074
rect 10108 13020 10164 13022
rect 9212 11394 9268 11396
rect 9212 11342 9214 11394
rect 9214 11342 9266 11394
rect 9266 11342 9268 11394
rect 9212 11340 9268 11342
rect 8764 11004 8820 11060
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 9100 10722 9156 10724
rect 9100 10670 9102 10722
rect 9102 10670 9154 10722
rect 9154 10670 9156 10722
rect 9100 10668 9156 10670
rect 9436 9938 9492 9940
rect 9436 9886 9438 9938
rect 9438 9886 9490 9938
rect 9490 9886 9492 9938
rect 9436 9884 9492 9886
rect 8988 9714 9044 9716
rect 8988 9662 8990 9714
rect 8990 9662 9042 9714
rect 9042 9662 9044 9714
rect 8988 9660 9044 9662
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 9772 11394 9828 11396
rect 9772 11342 9774 11394
rect 9774 11342 9826 11394
rect 9826 11342 9828 11394
rect 9772 11340 9828 11342
rect 10220 12290 10276 12292
rect 10220 12238 10222 12290
rect 10222 12238 10274 12290
rect 10274 12238 10276 12290
rect 10220 12236 10276 12238
rect 11004 18620 11060 18676
rect 11004 18172 11060 18228
rect 11564 20076 11620 20132
rect 11452 19964 11508 20020
rect 11340 19906 11396 19908
rect 11340 19854 11342 19906
rect 11342 19854 11394 19906
rect 11394 19854 11396 19906
rect 11340 19852 11396 19854
rect 11340 18674 11396 18676
rect 11340 18622 11342 18674
rect 11342 18622 11394 18674
rect 11394 18622 11396 18674
rect 11340 18620 11396 18622
rect 11452 18508 11508 18564
rect 11340 18172 11396 18228
rect 11340 17724 11396 17780
rect 10556 14700 10612 14756
rect 10892 14418 10948 14420
rect 10892 14366 10894 14418
rect 10894 14366 10946 14418
rect 10946 14366 10948 14418
rect 10892 14364 10948 14366
rect 11116 17052 11172 17108
rect 11004 13634 11060 13636
rect 11004 13582 11006 13634
rect 11006 13582 11058 13634
rect 11058 13582 11060 13634
rect 11004 13580 11060 13582
rect 10892 13468 10948 13524
rect 11228 16604 11284 16660
rect 11788 21196 11844 21252
rect 11788 20802 11844 20804
rect 11788 20750 11790 20802
rect 11790 20750 11842 20802
rect 11842 20750 11844 20802
rect 11788 20748 11844 20750
rect 12012 20972 12068 21028
rect 11900 20300 11956 20356
rect 12012 20076 12068 20132
rect 12012 19234 12068 19236
rect 12012 19182 12014 19234
rect 12014 19182 12066 19234
rect 12066 19182 12068 19234
rect 12012 19180 12068 19182
rect 12236 25506 12292 25508
rect 12236 25454 12238 25506
rect 12238 25454 12290 25506
rect 12290 25454 12292 25506
rect 12236 25452 12292 25454
rect 12460 25394 12516 25396
rect 12460 25342 12462 25394
rect 12462 25342 12514 25394
rect 12514 25342 12516 25394
rect 12460 25340 12516 25342
rect 13244 27244 13300 27300
rect 13804 27244 13860 27300
rect 13020 26124 13076 26180
rect 13356 26908 13412 26964
rect 12684 25506 12740 25508
rect 12684 25454 12686 25506
rect 12686 25454 12738 25506
rect 12738 25454 12740 25506
rect 12684 25452 12740 25454
rect 13020 25394 13076 25396
rect 13020 25342 13022 25394
rect 13022 25342 13074 25394
rect 13074 25342 13076 25394
rect 13020 25340 13076 25342
rect 12908 24892 12964 24948
rect 12684 24444 12740 24500
rect 12236 22428 12292 22484
rect 12460 22370 12516 22372
rect 12460 22318 12462 22370
rect 12462 22318 12514 22370
rect 12514 22318 12516 22370
rect 12460 22316 12516 22318
rect 12348 21868 12404 21924
rect 12236 21084 12292 21140
rect 12236 20636 12292 20692
rect 12236 19068 12292 19124
rect 11676 18844 11732 18900
rect 11564 17052 11620 17108
rect 11676 17724 11732 17780
rect 11452 15484 11508 15540
rect 11788 15484 11844 15540
rect 12348 16380 12404 16436
rect 12572 21196 12628 21252
rect 13020 24834 13076 24836
rect 13020 24782 13022 24834
rect 13022 24782 13074 24834
rect 13074 24782 13076 24834
rect 13020 24780 13076 24782
rect 12908 24220 12964 24276
rect 13468 26460 13524 26516
rect 13692 26962 13748 26964
rect 13692 26910 13694 26962
rect 13694 26910 13746 26962
rect 13746 26910 13748 26962
rect 13692 26908 13748 26910
rect 13580 26236 13636 26292
rect 14028 27804 14084 27860
rect 14028 27468 14084 27524
rect 13916 26684 13972 26740
rect 13916 26460 13972 26516
rect 13468 26178 13524 26180
rect 13468 26126 13470 26178
rect 13470 26126 13522 26178
rect 13522 26126 13524 26178
rect 13468 26124 13524 26126
rect 13692 25900 13748 25956
rect 13804 25564 13860 25620
rect 13916 25506 13972 25508
rect 13916 25454 13918 25506
rect 13918 25454 13970 25506
rect 13970 25454 13972 25506
rect 13916 25452 13972 25454
rect 13580 25004 13636 25060
rect 13468 24892 13524 24948
rect 13356 24220 13412 24276
rect 13468 21868 13524 21924
rect 13132 21532 13188 21588
rect 12684 21084 12740 21140
rect 11788 15036 11844 15092
rect 11228 13916 11284 13972
rect 10780 12066 10836 12068
rect 10780 12014 10782 12066
rect 10782 12014 10834 12066
rect 10834 12014 10836 12066
rect 10780 12012 10836 12014
rect 10444 11676 10500 11732
rect 10108 11116 10164 11172
rect 10220 11340 10276 11396
rect 10556 10892 10612 10948
rect 10444 10780 10500 10836
rect 10556 10498 10612 10500
rect 10556 10446 10558 10498
rect 10558 10446 10610 10498
rect 10610 10446 10612 10498
rect 10556 10444 10612 10446
rect 10332 9826 10388 9828
rect 10332 9774 10334 9826
rect 10334 9774 10386 9826
rect 10386 9774 10388 9826
rect 10332 9772 10388 9774
rect 9996 9324 10052 9380
rect 11788 13916 11844 13972
rect 11340 13746 11396 13748
rect 11340 13694 11342 13746
rect 11342 13694 11394 13746
rect 11394 13694 11396 13746
rect 11340 13692 11396 13694
rect 11228 12348 11284 12404
rect 11340 12124 11396 12180
rect 11228 11564 11284 11620
rect 11116 9324 11172 9380
rect 10892 9266 10948 9268
rect 10892 9214 10894 9266
rect 10894 9214 10946 9266
rect 10946 9214 10948 9266
rect 10892 9212 10948 9214
rect 10444 9042 10500 9044
rect 10444 8990 10446 9042
rect 10446 8990 10498 9042
rect 10498 8990 10500 9042
rect 10444 8988 10500 8990
rect 9884 8204 9940 8260
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 11004 7474 11060 7476
rect 11004 7422 11006 7474
rect 11006 7422 11058 7474
rect 11058 7422 11060 7474
rect 11004 7420 11060 7422
rect 10892 6972 10948 7028
rect 9884 6802 9940 6804
rect 9884 6750 9886 6802
rect 9886 6750 9938 6802
rect 9938 6750 9940 6802
rect 9884 6748 9940 6750
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 11452 10610 11508 10612
rect 11452 10558 11454 10610
rect 11454 10558 11506 10610
rect 11506 10558 11508 10610
rect 11452 10556 11508 10558
rect 11900 13692 11956 13748
rect 12124 14364 12180 14420
rect 12012 12460 12068 12516
rect 12684 20188 12740 20244
rect 12908 19964 12964 20020
rect 12796 19852 12852 19908
rect 12572 19740 12628 19796
rect 12572 18956 12628 19012
rect 13020 18844 13076 18900
rect 13916 24108 13972 24164
rect 13916 23714 13972 23716
rect 13916 23662 13918 23714
rect 13918 23662 13970 23714
rect 13970 23662 13972 23714
rect 13916 23660 13972 23662
rect 13916 23324 13972 23380
rect 13692 21532 13748 21588
rect 13804 22540 13860 22596
rect 13132 18396 13188 18452
rect 13356 21420 13412 21476
rect 13468 20690 13524 20692
rect 13468 20638 13470 20690
rect 13470 20638 13522 20690
rect 13522 20638 13524 20690
rect 13468 20636 13524 20638
rect 13692 20524 13748 20580
rect 13916 22204 13972 22260
rect 13356 18844 13412 18900
rect 13468 19516 13524 19572
rect 13692 20018 13748 20020
rect 13692 19966 13694 20018
rect 13694 19966 13746 20018
rect 13746 19966 13748 20018
rect 13692 19964 13748 19966
rect 13916 19740 13972 19796
rect 13468 18620 13524 18676
rect 13692 18450 13748 18452
rect 13692 18398 13694 18450
rect 13694 18398 13746 18450
rect 13746 18398 13748 18450
rect 13692 18396 13748 18398
rect 13580 18284 13636 18340
rect 12908 17554 12964 17556
rect 12908 17502 12910 17554
rect 12910 17502 12962 17554
rect 12962 17502 12964 17554
rect 12908 17500 12964 17502
rect 14364 29426 14420 29428
rect 14364 29374 14366 29426
rect 14366 29374 14418 29426
rect 14418 29374 14420 29426
rect 14364 29372 14420 29374
rect 15372 29372 15428 29428
rect 14700 28642 14756 28644
rect 14700 28590 14702 28642
rect 14702 28590 14754 28642
rect 14754 28590 14756 28642
rect 14700 28588 14756 28590
rect 14364 27746 14420 27748
rect 14364 27694 14366 27746
rect 14366 27694 14418 27746
rect 14418 27694 14420 27746
rect 14364 27692 14420 27694
rect 15596 29426 15652 29428
rect 15596 29374 15598 29426
rect 15598 29374 15650 29426
rect 15650 29374 15652 29426
rect 15596 29372 15652 29374
rect 15484 28642 15540 28644
rect 15484 28590 15486 28642
rect 15486 28590 15538 28642
rect 15538 28590 15540 28642
rect 15484 28588 15540 28590
rect 16716 29314 16772 29316
rect 16716 29262 16718 29314
rect 16718 29262 16770 29314
rect 16770 29262 16772 29314
rect 16716 29260 16772 29262
rect 16044 28700 16100 28756
rect 16380 28700 16436 28756
rect 15596 28476 15652 28532
rect 15148 27916 15204 27972
rect 14252 27132 14308 27188
rect 14252 26684 14308 26740
rect 14252 26012 14308 26068
rect 14140 25788 14196 25844
rect 14700 27132 14756 27188
rect 14364 25564 14420 25620
rect 14476 25676 14532 25732
rect 14140 24892 14196 24948
rect 14252 25452 14308 25508
rect 14252 23324 14308 23380
rect 14364 24610 14420 24612
rect 14364 24558 14366 24610
rect 14366 24558 14418 24610
rect 14418 24558 14420 24610
rect 14364 24556 14420 24558
rect 15708 27074 15764 27076
rect 15708 27022 15710 27074
rect 15710 27022 15762 27074
rect 15762 27022 15764 27074
rect 15708 27020 15764 27022
rect 16716 28530 16772 28532
rect 16716 28478 16718 28530
rect 16718 28478 16770 28530
rect 16770 28478 16772 28530
rect 16716 28476 16772 28478
rect 16268 27970 16324 27972
rect 16268 27918 16270 27970
rect 16270 27918 16322 27970
rect 16322 27918 16324 27970
rect 16268 27916 16324 27918
rect 16268 27298 16324 27300
rect 16268 27246 16270 27298
rect 16270 27246 16322 27298
rect 16322 27246 16324 27298
rect 16268 27244 16324 27246
rect 15372 26572 15428 26628
rect 15260 26290 15316 26292
rect 15260 26238 15262 26290
rect 15262 26238 15314 26290
rect 15314 26238 15316 26290
rect 15260 26236 15316 26238
rect 14812 25900 14868 25956
rect 14812 25564 14868 25620
rect 14812 25116 14868 25172
rect 14700 25004 14756 25060
rect 14140 21644 14196 21700
rect 14140 20636 14196 20692
rect 14252 19234 14308 19236
rect 14252 19182 14254 19234
rect 14254 19182 14306 19234
rect 14306 19182 14308 19234
rect 14252 19180 14308 19182
rect 14028 19068 14084 19124
rect 15596 26012 15652 26068
rect 15372 25900 15428 25956
rect 15372 25452 15428 25508
rect 15036 25116 15092 25172
rect 16268 26908 16324 26964
rect 16156 26290 16212 26292
rect 16156 26238 16158 26290
rect 16158 26238 16210 26290
rect 16210 26238 16212 26290
rect 16156 26236 16212 26238
rect 16268 25788 16324 25844
rect 15932 25506 15988 25508
rect 15932 25454 15934 25506
rect 15934 25454 15986 25506
rect 15986 25454 15988 25506
rect 15932 25452 15988 25454
rect 15820 25116 15876 25172
rect 14924 24220 14980 24276
rect 15708 25004 15764 25060
rect 14700 23772 14756 23828
rect 14588 20860 14644 20916
rect 14476 19964 14532 20020
rect 14476 19292 14532 19348
rect 13580 16828 13636 16884
rect 13468 16770 13524 16772
rect 13468 16718 13470 16770
rect 13470 16718 13522 16770
rect 13522 16718 13524 16770
rect 13468 16716 13524 16718
rect 13356 16156 13412 16212
rect 13692 16492 13748 16548
rect 13580 16098 13636 16100
rect 13580 16046 13582 16098
rect 13582 16046 13634 16098
rect 13634 16046 13636 16098
rect 13580 16044 13636 16046
rect 12572 15708 12628 15764
rect 13580 15708 13636 15764
rect 13132 15484 13188 15540
rect 12908 14924 12964 14980
rect 12572 14530 12628 14532
rect 12572 14478 12574 14530
rect 12574 14478 12626 14530
rect 12626 14478 12628 14530
rect 12572 14476 12628 14478
rect 12684 14364 12740 14420
rect 13692 15260 13748 15316
rect 13468 14588 13524 14644
rect 11900 12236 11956 12292
rect 12348 12796 12404 12852
rect 11676 12124 11732 12180
rect 11340 8930 11396 8932
rect 11340 8878 11342 8930
rect 11342 8878 11394 8930
rect 11394 8878 11396 8930
rect 11340 8876 11396 8878
rect 11340 8652 11396 8708
rect 11676 9996 11732 10052
rect 11900 11564 11956 11620
rect 11900 11394 11956 11396
rect 11900 11342 11902 11394
rect 11902 11342 11954 11394
rect 11954 11342 11956 11394
rect 11900 11340 11956 11342
rect 12348 11282 12404 11284
rect 12348 11230 12350 11282
rect 12350 11230 12402 11282
rect 12402 11230 12404 11282
rect 12348 11228 12404 11230
rect 12348 10556 12404 10612
rect 12908 13074 12964 13076
rect 12908 13022 12910 13074
rect 12910 13022 12962 13074
rect 12962 13022 12964 13074
rect 12908 13020 12964 13022
rect 12796 11676 12852 11732
rect 12908 11116 12964 11172
rect 12572 10780 12628 10836
rect 12236 9826 12292 9828
rect 12236 9774 12238 9826
rect 12238 9774 12290 9826
rect 12290 9774 12292 9826
rect 12236 9772 12292 9774
rect 11676 8876 11732 8932
rect 11676 7420 11732 7476
rect 11340 6578 11396 6580
rect 11340 6526 11342 6578
rect 11342 6526 11394 6578
rect 11394 6526 11396 6578
rect 11340 6524 11396 6526
rect 4732 3276 4788 3332
rect 5516 3330 5572 3332
rect 5516 3278 5518 3330
rect 5518 3278 5570 3330
rect 5570 3278 5572 3330
rect 5516 3276 5572 3278
rect 11564 3276 11620 3332
rect 12012 8092 12068 8148
rect 12236 8876 12292 8932
rect 12796 10892 12852 10948
rect 12908 10780 12964 10836
rect 12796 9884 12852 9940
rect 12684 8930 12740 8932
rect 12684 8878 12686 8930
rect 12686 8878 12738 8930
rect 12738 8878 12740 8930
rect 12684 8876 12740 8878
rect 12348 8652 12404 8708
rect 13020 8540 13076 8596
rect 13244 13020 13300 13076
rect 13692 14812 13748 14868
rect 13692 14028 13748 14084
rect 13692 12738 13748 12740
rect 13692 12686 13694 12738
rect 13694 12686 13746 12738
rect 13746 12686 13748 12738
rect 13692 12684 13748 12686
rect 13916 16828 13972 16884
rect 14028 15874 14084 15876
rect 14028 15822 14030 15874
rect 14030 15822 14082 15874
rect 14082 15822 14084 15874
rect 14028 15820 14084 15822
rect 14140 15596 14196 15652
rect 16268 24892 16324 24948
rect 15932 24220 15988 24276
rect 14812 20076 14868 20132
rect 15708 23884 15764 23940
rect 16044 23996 16100 24052
rect 15372 21308 15428 21364
rect 15036 20860 15092 20916
rect 16268 23436 16324 23492
rect 16156 23042 16212 23044
rect 16156 22990 16158 23042
rect 16158 22990 16210 23042
rect 16210 22990 16212 23042
rect 16156 22988 16212 22990
rect 16828 27356 16884 27412
rect 16604 27186 16660 27188
rect 16604 27134 16606 27186
rect 16606 27134 16658 27186
rect 16658 27134 16660 27186
rect 16604 27132 16660 27134
rect 16716 26236 16772 26292
rect 16492 25228 16548 25284
rect 16604 24610 16660 24612
rect 16604 24558 16606 24610
rect 16606 24558 16658 24610
rect 16658 24558 16660 24610
rect 16604 24556 16660 24558
rect 16828 26178 16884 26180
rect 16828 26126 16830 26178
rect 16830 26126 16882 26178
rect 16882 26126 16884 26178
rect 16828 26124 16884 26126
rect 17500 29484 17556 29540
rect 17724 29596 17780 29652
rect 17612 29426 17668 29428
rect 17612 29374 17614 29426
rect 17614 29374 17666 29426
rect 17666 29374 17668 29426
rect 17612 29372 17668 29374
rect 19180 32844 19236 32900
rect 18956 31164 19012 31220
rect 19180 31164 19236 31220
rect 21644 45724 21700 45780
rect 21532 45388 21588 45444
rect 22428 53618 22484 53620
rect 22428 53566 22430 53618
rect 22430 53566 22482 53618
rect 22482 53566 22484 53618
rect 22428 53564 22484 53566
rect 22540 53058 22596 53060
rect 22540 53006 22542 53058
rect 22542 53006 22594 53058
rect 22594 53006 22596 53058
rect 22540 53004 22596 53006
rect 22540 52162 22596 52164
rect 22540 52110 22542 52162
rect 22542 52110 22594 52162
rect 22594 52110 22596 52162
rect 22540 52108 22596 52110
rect 24780 56364 24836 56420
rect 23324 56306 23380 56308
rect 23324 56254 23326 56306
rect 23326 56254 23378 56306
rect 23378 56254 23380 56306
rect 23324 56252 23380 56254
rect 24668 56194 24724 56196
rect 24668 56142 24670 56194
rect 24670 56142 24722 56194
rect 24722 56142 24724 56194
rect 24668 56140 24724 56142
rect 23548 56028 23604 56084
rect 23212 55468 23268 55524
rect 23100 53788 23156 53844
rect 22988 53564 23044 53620
rect 24556 55804 24612 55860
rect 24332 55410 24388 55412
rect 24332 55358 24334 55410
rect 24334 55358 24386 55410
rect 24386 55358 24388 55410
rect 24332 55356 24388 55358
rect 23548 55132 23604 55188
rect 23772 54796 23828 54852
rect 23548 54348 23604 54404
rect 23436 53788 23492 53844
rect 22988 52220 23044 52276
rect 22316 51436 22372 51492
rect 22204 50540 22260 50596
rect 22540 51154 22596 51156
rect 22540 51102 22542 51154
rect 22542 51102 22594 51154
rect 22594 51102 22596 51154
rect 22540 51100 22596 51102
rect 22092 49644 22148 49700
rect 21868 48076 21924 48132
rect 22316 47628 22372 47684
rect 21868 46956 21924 47012
rect 21868 46172 21924 46228
rect 22092 46060 22148 46116
rect 21644 43426 21700 43428
rect 21644 43374 21646 43426
rect 21646 43374 21698 43426
rect 21698 43374 21700 43426
rect 21644 43372 21700 43374
rect 21420 43260 21476 43316
rect 21868 44322 21924 44324
rect 21868 44270 21870 44322
rect 21870 44270 21922 44322
rect 21922 44270 21924 44322
rect 21868 44268 21924 44270
rect 21756 43260 21812 43316
rect 21868 44044 21924 44100
rect 21980 43148 22036 43204
rect 23324 52780 23380 52836
rect 23548 53340 23604 53396
rect 22876 51378 22932 51380
rect 22876 51326 22878 51378
rect 22878 51326 22930 51378
rect 22930 51326 22932 51378
rect 22876 51324 22932 51326
rect 22988 50316 23044 50372
rect 22988 49980 23044 50036
rect 22764 49810 22820 49812
rect 22764 49758 22766 49810
rect 22766 49758 22818 49810
rect 22818 49758 22820 49810
rect 22764 49756 22820 49758
rect 23100 49868 23156 49924
rect 23884 54348 23940 54404
rect 23660 52556 23716 52612
rect 23548 51324 23604 51380
rect 23660 52108 23716 52164
rect 23324 49420 23380 49476
rect 23548 51100 23604 51156
rect 23324 48972 23380 49028
rect 22764 48748 22820 48804
rect 22764 47458 22820 47460
rect 22764 47406 22766 47458
rect 22766 47406 22818 47458
rect 22818 47406 22820 47458
rect 22764 47404 22820 47406
rect 22876 48636 22932 48692
rect 24556 54514 24612 54516
rect 24556 54462 24558 54514
rect 24558 54462 24610 54514
rect 24610 54462 24612 54514
rect 24556 54460 24612 54462
rect 24780 55804 24836 55860
rect 24668 54348 24724 54404
rect 24220 54290 24276 54292
rect 24220 54238 24222 54290
rect 24222 54238 24274 54290
rect 24274 54238 24276 54290
rect 24220 54236 24276 54238
rect 24108 53730 24164 53732
rect 24108 53678 24110 53730
rect 24110 53678 24162 53730
rect 24162 53678 24164 53730
rect 24108 53676 24164 53678
rect 23996 52108 24052 52164
rect 24668 53452 24724 53508
rect 24332 53170 24388 53172
rect 24332 53118 24334 53170
rect 24334 53118 24386 53170
rect 24386 53118 24388 53170
rect 24332 53116 24388 53118
rect 24444 53004 24500 53060
rect 24892 54796 24948 54852
rect 24668 53058 24724 53060
rect 24668 53006 24670 53058
rect 24670 53006 24722 53058
rect 24722 53006 24724 53058
rect 24668 53004 24724 53006
rect 24108 51660 24164 51716
rect 23884 50764 23940 50820
rect 23772 50652 23828 50708
rect 24780 52556 24836 52612
rect 24220 51378 24276 51380
rect 24220 51326 24222 51378
rect 24222 51326 24274 51378
rect 24274 51326 24276 51378
rect 24220 51324 24276 51326
rect 23996 50540 24052 50596
rect 24108 51212 24164 51268
rect 24332 50594 24388 50596
rect 24332 50542 24334 50594
rect 24334 50542 24386 50594
rect 24386 50542 24388 50594
rect 24332 50540 24388 50542
rect 24444 50428 24500 50484
rect 23660 49922 23716 49924
rect 23660 49870 23662 49922
rect 23662 49870 23714 49922
rect 23714 49870 23716 49922
rect 23660 49868 23716 49870
rect 22540 47068 22596 47124
rect 22428 45836 22484 45892
rect 22204 45500 22260 45556
rect 21532 42866 21588 42868
rect 21532 42814 21534 42866
rect 21534 42814 21586 42866
rect 21586 42814 21588 42866
rect 21532 42812 21588 42814
rect 21308 42028 21364 42084
rect 21532 42476 21588 42532
rect 21084 41580 21140 41636
rect 21196 41020 21252 41076
rect 21756 42140 21812 42196
rect 23100 48076 23156 48132
rect 22988 47404 23044 47460
rect 22764 46060 22820 46116
rect 22652 45164 22708 45220
rect 22764 45612 22820 45668
rect 22316 43596 22372 43652
rect 22316 43372 22372 43428
rect 22092 42588 22148 42644
rect 22764 43426 22820 43428
rect 22764 43374 22766 43426
rect 22766 43374 22818 43426
rect 22818 43374 22820 43426
rect 22764 43372 22820 43374
rect 23100 47292 23156 47348
rect 23212 47068 23268 47124
rect 22988 44268 23044 44324
rect 22316 42028 22372 42084
rect 22428 41916 22484 41972
rect 22092 41580 22148 41636
rect 22316 41356 22372 41412
rect 21756 41244 21812 41300
rect 22540 41298 22596 41300
rect 22540 41246 22542 41298
rect 22542 41246 22594 41298
rect 22594 41246 22596 41298
rect 22540 41244 22596 41246
rect 22652 41692 22708 41748
rect 22092 41020 22148 41076
rect 21196 40514 21252 40516
rect 21196 40462 21198 40514
rect 21198 40462 21250 40514
rect 21250 40462 21252 40514
rect 21196 40460 21252 40462
rect 21644 40796 21700 40852
rect 21308 40236 21364 40292
rect 21084 39004 21140 39060
rect 21084 38108 21140 38164
rect 21308 37826 21364 37828
rect 21308 37774 21310 37826
rect 21310 37774 21362 37826
rect 21362 37774 21364 37826
rect 21308 37772 21364 37774
rect 22204 40626 22260 40628
rect 22204 40574 22206 40626
rect 22206 40574 22258 40626
rect 22258 40574 22260 40626
rect 22204 40572 22260 40574
rect 21644 40012 21700 40068
rect 23100 44098 23156 44100
rect 23100 44046 23102 44098
rect 23102 44046 23154 44098
rect 23154 44046 23156 44098
rect 23100 44044 23156 44046
rect 23212 43372 23268 43428
rect 22876 41468 22932 41524
rect 23100 41356 23156 41412
rect 24108 49308 24164 49364
rect 24220 48972 24276 49028
rect 24668 49922 24724 49924
rect 24668 49870 24670 49922
rect 24670 49870 24722 49922
rect 24722 49870 24724 49922
rect 24668 49868 24724 49870
rect 24556 49308 24612 49364
rect 24332 48748 24388 48804
rect 24892 50876 24948 50932
rect 26460 57148 26516 57204
rect 25564 56194 25620 56196
rect 25564 56142 25566 56194
rect 25566 56142 25618 56194
rect 25618 56142 25620 56194
rect 25564 56140 25620 56142
rect 25228 55916 25284 55972
rect 26124 55356 26180 55412
rect 25340 55244 25396 55300
rect 26236 54738 26292 54740
rect 26236 54686 26238 54738
rect 26238 54686 26290 54738
rect 26290 54686 26292 54738
rect 26236 54684 26292 54686
rect 26124 54348 26180 54404
rect 26012 53676 26068 53732
rect 25116 53004 25172 53060
rect 24892 50706 24948 50708
rect 24892 50654 24894 50706
rect 24894 50654 24946 50706
rect 24946 50654 24948 50706
rect 24892 50652 24948 50654
rect 24220 48466 24276 48468
rect 24220 48414 24222 48466
rect 24222 48414 24274 48466
rect 24274 48414 24276 48466
rect 24220 48412 24276 48414
rect 23772 47458 23828 47460
rect 23772 47406 23774 47458
rect 23774 47406 23826 47458
rect 23826 47406 23828 47458
rect 23772 47404 23828 47406
rect 24108 48076 24164 48132
rect 24108 47516 24164 47572
rect 23996 46732 24052 46788
rect 23772 46674 23828 46676
rect 23772 46622 23774 46674
rect 23774 46622 23826 46674
rect 23826 46622 23828 46674
rect 23772 46620 23828 46622
rect 23884 46284 23940 46340
rect 23884 46002 23940 46004
rect 23884 45950 23886 46002
rect 23886 45950 23938 46002
rect 23938 45950 23940 46002
rect 23884 45948 23940 45950
rect 23660 45724 23716 45780
rect 23436 45666 23492 45668
rect 23436 45614 23438 45666
rect 23438 45614 23490 45666
rect 23490 45614 23492 45666
rect 23436 45612 23492 45614
rect 23436 44492 23492 44548
rect 23996 45388 24052 45444
rect 23772 44380 23828 44436
rect 23548 44098 23604 44100
rect 23548 44046 23550 44098
rect 23550 44046 23602 44098
rect 23602 44046 23604 44098
rect 23548 44044 23604 44046
rect 23884 44604 23940 44660
rect 24108 44322 24164 44324
rect 24108 44270 24110 44322
rect 24110 44270 24162 44322
rect 24162 44270 24164 44322
rect 24108 44268 24164 44270
rect 23436 43650 23492 43652
rect 23436 43598 23438 43650
rect 23438 43598 23490 43650
rect 23490 43598 23492 43650
rect 23436 43596 23492 43598
rect 23548 42700 23604 42756
rect 23436 41468 23492 41524
rect 23436 40908 23492 40964
rect 22652 40460 22708 40516
rect 22428 40012 22484 40068
rect 22652 39842 22708 39844
rect 22652 39790 22654 39842
rect 22654 39790 22706 39842
rect 22706 39790 22708 39842
rect 22652 39788 22708 39790
rect 22428 39730 22484 39732
rect 22428 39678 22430 39730
rect 22430 39678 22482 39730
rect 22482 39678 22484 39730
rect 22428 39676 22484 39678
rect 22092 39618 22148 39620
rect 22092 39566 22094 39618
rect 22094 39566 22146 39618
rect 22146 39566 22148 39618
rect 22092 39564 22148 39566
rect 22204 39340 22260 39396
rect 23100 39730 23156 39732
rect 23100 39678 23102 39730
rect 23102 39678 23154 39730
rect 23154 39678 23156 39730
rect 23100 39676 23156 39678
rect 22652 39340 22708 39396
rect 22316 38780 22372 38836
rect 22204 38556 22260 38612
rect 21868 37660 21924 37716
rect 22092 37884 22148 37940
rect 20972 37212 21028 37268
rect 20748 36594 20804 36596
rect 20748 36542 20750 36594
rect 20750 36542 20802 36594
rect 20802 36542 20804 36594
rect 20748 36540 20804 36542
rect 20636 34748 20692 34804
rect 20636 34412 20692 34468
rect 19516 33740 19572 33796
rect 19516 33570 19572 33572
rect 19516 33518 19518 33570
rect 19518 33518 19570 33570
rect 19570 33518 19572 33570
rect 19516 33516 19572 33518
rect 20524 33852 20580 33908
rect 20412 33292 20468 33348
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19852 32674 19908 32676
rect 19852 32622 19854 32674
rect 19854 32622 19906 32674
rect 19906 32622 19908 32674
rect 19852 32620 19908 32622
rect 18956 30994 19012 30996
rect 18956 30942 18958 30994
rect 18958 30942 19010 30994
rect 19010 30942 19012 30994
rect 18956 30940 19012 30942
rect 19180 30380 19236 30436
rect 17948 29538 18004 29540
rect 17948 29486 17950 29538
rect 17950 29486 18002 29538
rect 18002 29486 18004 29538
rect 17948 29484 18004 29486
rect 17836 29426 17892 29428
rect 17836 29374 17838 29426
rect 17838 29374 17890 29426
rect 17890 29374 17892 29426
rect 17836 29372 17892 29374
rect 18060 29372 18116 29428
rect 19964 31500 20020 31556
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19404 30994 19460 30996
rect 19404 30942 19406 30994
rect 19406 30942 19458 30994
rect 19458 30942 19460 30994
rect 19404 30940 19460 30942
rect 20076 30380 20132 30436
rect 19404 30210 19460 30212
rect 19404 30158 19406 30210
rect 19406 30158 19458 30210
rect 19458 30158 19460 30210
rect 19404 30156 19460 30158
rect 19292 30044 19348 30100
rect 20076 30210 20132 30212
rect 20076 30158 20078 30210
rect 20078 30158 20130 30210
rect 20130 30158 20132 30210
rect 20076 30156 20132 30158
rect 20860 33292 20916 33348
rect 21868 37266 21924 37268
rect 21868 37214 21870 37266
rect 21870 37214 21922 37266
rect 21922 37214 21924 37266
rect 21868 37212 21924 37214
rect 21308 36652 21364 36708
rect 21420 36876 21476 36932
rect 22092 36876 22148 36932
rect 21532 36594 21588 36596
rect 21532 36542 21534 36594
rect 21534 36542 21586 36594
rect 21586 36542 21588 36594
rect 21532 36540 21588 36542
rect 21420 36316 21476 36372
rect 22316 38108 22372 38164
rect 22876 37996 22932 38052
rect 22988 37884 23044 37940
rect 22988 37548 23044 37604
rect 22316 36540 22372 36596
rect 21308 35644 21364 35700
rect 22764 35810 22820 35812
rect 22764 35758 22766 35810
rect 22766 35758 22818 35810
rect 22818 35758 22820 35810
rect 22764 35756 22820 35758
rect 23324 40012 23380 40068
rect 23324 39228 23380 39284
rect 23660 42082 23716 42084
rect 23660 42030 23662 42082
rect 23662 42030 23714 42082
rect 23714 42030 23716 42082
rect 23660 42028 23716 42030
rect 23884 43484 23940 43540
rect 23884 43148 23940 43204
rect 24668 48354 24724 48356
rect 24668 48302 24670 48354
rect 24670 48302 24722 48354
rect 24722 48302 24724 48354
rect 24668 48300 24724 48302
rect 24444 45778 24500 45780
rect 24444 45726 24446 45778
rect 24446 45726 24498 45778
rect 24498 45726 24500 45778
rect 24444 45724 24500 45726
rect 24444 45218 24500 45220
rect 24444 45166 24446 45218
rect 24446 45166 24498 45218
rect 24498 45166 24500 45218
rect 24444 45164 24500 45166
rect 24668 47570 24724 47572
rect 24668 47518 24670 47570
rect 24670 47518 24722 47570
rect 24722 47518 24724 47570
rect 24668 47516 24724 47518
rect 25564 52834 25620 52836
rect 25564 52782 25566 52834
rect 25566 52782 25618 52834
rect 25618 52782 25620 52834
rect 25564 52780 25620 52782
rect 25228 51602 25284 51604
rect 25228 51550 25230 51602
rect 25230 51550 25282 51602
rect 25282 51550 25284 51602
rect 25228 51548 25284 51550
rect 25228 51324 25284 51380
rect 26012 52332 26068 52388
rect 25676 52108 25732 52164
rect 25564 50540 25620 50596
rect 26124 51996 26180 52052
rect 26124 51378 26180 51380
rect 26124 51326 26126 51378
rect 26126 51326 26178 51378
rect 26178 51326 26180 51378
rect 26124 51324 26180 51326
rect 26124 50764 26180 50820
rect 25788 50652 25844 50708
rect 25900 50204 25956 50260
rect 25676 50092 25732 50148
rect 26012 50092 26068 50148
rect 25564 49868 25620 49924
rect 26012 49420 26068 49476
rect 26012 48972 26068 49028
rect 25676 48860 25732 48916
rect 25900 48748 25956 48804
rect 25564 48188 25620 48244
rect 25340 47852 25396 47908
rect 25228 47404 25284 47460
rect 25788 47964 25844 48020
rect 25676 47852 25732 47908
rect 25676 47628 25732 47684
rect 25452 47292 25508 47348
rect 24668 46284 24724 46340
rect 24892 46620 24948 46676
rect 24780 46060 24836 46116
rect 24668 45388 24724 45444
rect 24780 45218 24836 45220
rect 24780 45166 24782 45218
rect 24782 45166 24834 45218
rect 24834 45166 24836 45218
rect 24780 45164 24836 45166
rect 24556 44492 24612 44548
rect 25228 46060 25284 46116
rect 26236 50316 26292 50372
rect 26012 47458 26068 47460
rect 26012 47406 26014 47458
rect 26014 47406 26066 47458
rect 26066 47406 26068 47458
rect 26012 47404 26068 47406
rect 25564 46508 25620 46564
rect 25340 45612 25396 45668
rect 25340 45388 25396 45444
rect 25452 45164 25508 45220
rect 25116 45052 25172 45108
rect 24892 44380 24948 44436
rect 25228 44604 25284 44660
rect 24332 43650 24388 43652
rect 24332 43598 24334 43650
rect 24334 43598 24386 43650
rect 24386 43598 24388 43650
rect 24332 43596 24388 43598
rect 24556 44322 24612 44324
rect 24556 44270 24558 44322
rect 24558 44270 24610 44322
rect 24610 44270 24612 44322
rect 24556 44268 24612 44270
rect 24108 43148 24164 43204
rect 23884 42700 23940 42756
rect 24444 42754 24500 42756
rect 24444 42702 24446 42754
rect 24446 42702 24498 42754
rect 24498 42702 24500 42754
rect 24444 42700 24500 42702
rect 24108 42364 24164 42420
rect 23772 38892 23828 38948
rect 24220 41580 24276 41636
rect 25004 44322 25060 44324
rect 25004 44270 25006 44322
rect 25006 44270 25058 44322
rect 25058 44270 25060 44322
rect 25004 44268 25060 44270
rect 24892 43596 24948 43652
rect 24220 41020 24276 41076
rect 25340 44044 25396 44100
rect 25788 46172 25844 46228
rect 25676 45724 25732 45780
rect 25340 43538 25396 43540
rect 25340 43486 25342 43538
rect 25342 43486 25394 43538
rect 25394 43486 25396 43538
rect 25340 43484 25396 43486
rect 24780 40962 24836 40964
rect 24780 40910 24782 40962
rect 24782 40910 24834 40962
rect 24834 40910 24836 40962
rect 24780 40908 24836 40910
rect 24332 40402 24388 40404
rect 24332 40350 24334 40402
rect 24334 40350 24386 40402
rect 24386 40350 24388 40402
rect 24332 40348 24388 40350
rect 25004 40124 25060 40180
rect 23996 39340 24052 39396
rect 24220 39116 24276 39172
rect 24108 39004 24164 39060
rect 23884 38668 23940 38724
rect 23436 38050 23492 38052
rect 23436 37998 23438 38050
rect 23438 37998 23490 38050
rect 23490 37998 23492 38050
rect 23436 37996 23492 37998
rect 23772 38556 23828 38612
rect 23548 37772 23604 37828
rect 23548 37324 23604 37380
rect 23324 35980 23380 36036
rect 22428 35084 22484 35140
rect 21980 34972 22036 35028
rect 21308 34860 21364 34916
rect 22764 34972 22820 35028
rect 21532 34636 21588 34692
rect 21308 33852 21364 33908
rect 21420 34300 21476 34356
rect 21756 34354 21812 34356
rect 21756 34302 21758 34354
rect 21758 34302 21810 34354
rect 21810 34302 21812 34354
rect 21756 34300 21812 34302
rect 22988 34300 23044 34356
rect 21532 34130 21588 34132
rect 21532 34078 21534 34130
rect 21534 34078 21586 34130
rect 21586 34078 21588 34130
rect 21532 34076 21588 34078
rect 23548 35868 23604 35924
rect 23548 34412 23604 34468
rect 25116 39506 25172 39508
rect 25116 39454 25118 39506
rect 25118 39454 25170 39506
rect 25170 39454 25172 39506
rect 25116 39452 25172 39454
rect 25564 43036 25620 43092
rect 25788 43596 25844 43652
rect 30604 57596 30660 57652
rect 26684 57148 26740 57204
rect 27580 57260 27636 57316
rect 27020 56588 27076 56644
rect 26684 55356 26740 55412
rect 26796 54796 26852 54852
rect 26908 54514 26964 54516
rect 26908 54462 26910 54514
rect 26910 54462 26962 54514
rect 26962 54462 26964 54514
rect 26908 54460 26964 54462
rect 26460 53564 26516 53620
rect 26684 53730 26740 53732
rect 26684 53678 26686 53730
rect 26686 53678 26738 53730
rect 26738 53678 26740 53730
rect 26684 53676 26740 53678
rect 26572 53452 26628 53508
rect 26572 52834 26628 52836
rect 26572 52782 26574 52834
rect 26574 52782 26626 52834
rect 26626 52782 26628 52834
rect 26572 52780 26628 52782
rect 26460 52444 26516 52500
rect 27580 55244 27636 55300
rect 27580 55074 27636 55076
rect 27580 55022 27582 55074
rect 27582 55022 27634 55074
rect 27634 55022 27636 55074
rect 27580 55020 27636 55022
rect 27580 54124 27636 54180
rect 27916 55580 27972 55636
rect 28700 56194 28756 56196
rect 28700 56142 28702 56194
rect 28702 56142 28754 56194
rect 28754 56142 28756 56194
rect 28700 56140 28756 56142
rect 28700 55804 28756 55860
rect 28364 55468 28420 55524
rect 29484 55692 29540 55748
rect 26908 53452 26964 53508
rect 28252 55298 28308 55300
rect 28252 55246 28254 55298
rect 28254 55246 28306 55298
rect 28306 55246 28308 55298
rect 28252 55244 28308 55246
rect 28140 54012 28196 54068
rect 28140 53788 28196 53844
rect 28028 53506 28084 53508
rect 28028 53454 28030 53506
rect 28030 53454 28082 53506
rect 28082 53454 28084 53506
rect 28028 53452 28084 53454
rect 28364 54460 28420 54516
rect 28364 54236 28420 54292
rect 28364 53340 28420 53396
rect 28028 53116 28084 53172
rect 27356 52892 27412 52948
rect 26684 52332 26740 52388
rect 26796 52220 26852 52276
rect 26572 51266 26628 51268
rect 26572 51214 26574 51266
rect 26574 51214 26626 51266
rect 26626 51214 26628 51266
rect 26572 51212 26628 51214
rect 27132 52162 27188 52164
rect 27132 52110 27134 52162
rect 27134 52110 27186 52162
rect 27186 52110 27188 52162
rect 27132 52108 27188 52110
rect 27132 51378 27188 51380
rect 27132 51326 27134 51378
rect 27134 51326 27186 51378
rect 27186 51326 27188 51378
rect 27132 51324 27188 51326
rect 26460 50092 26516 50148
rect 26572 49922 26628 49924
rect 26572 49870 26574 49922
rect 26574 49870 26626 49922
rect 26626 49870 26628 49922
rect 26572 49868 26628 49870
rect 26348 47346 26404 47348
rect 26348 47294 26350 47346
rect 26350 47294 26402 47346
rect 26402 47294 26404 47346
rect 26348 47292 26404 47294
rect 26236 46620 26292 46676
rect 26572 48972 26628 49028
rect 27580 52556 27636 52612
rect 28028 52444 28084 52500
rect 27916 52220 27972 52276
rect 27804 51212 27860 51268
rect 26796 50316 26852 50372
rect 26908 50092 26964 50148
rect 26796 49756 26852 49812
rect 26796 49532 26852 49588
rect 26908 49308 26964 49364
rect 26684 48748 26740 48804
rect 26572 48412 26628 48468
rect 26572 47964 26628 48020
rect 26460 46620 26516 46676
rect 26796 48466 26852 48468
rect 26796 48414 26798 48466
rect 26798 48414 26850 48466
rect 26850 48414 26852 48466
rect 26796 48412 26852 48414
rect 26796 47852 26852 47908
rect 26684 46620 26740 46676
rect 26572 46562 26628 46564
rect 26572 46510 26574 46562
rect 26574 46510 26626 46562
rect 26626 46510 26628 46562
rect 26572 46508 26628 46510
rect 26236 46396 26292 46452
rect 26796 46396 26852 46452
rect 26572 45890 26628 45892
rect 26572 45838 26574 45890
rect 26574 45838 26626 45890
rect 26626 45838 26628 45890
rect 26572 45836 26628 45838
rect 26572 45388 26628 45444
rect 26236 44994 26292 44996
rect 26236 44942 26238 44994
rect 26238 44942 26290 44994
rect 26290 44942 26292 44994
rect 26236 44940 26292 44942
rect 26460 44156 26516 44212
rect 27356 50594 27412 50596
rect 27356 50542 27358 50594
rect 27358 50542 27410 50594
rect 27410 50542 27412 50594
rect 27356 50540 27412 50542
rect 27132 50316 27188 50372
rect 27356 50316 27412 50372
rect 27244 50092 27300 50148
rect 27468 50092 27524 50148
rect 27244 49810 27300 49812
rect 27244 49758 27246 49810
rect 27246 49758 27298 49810
rect 27298 49758 27300 49810
rect 27244 49756 27300 49758
rect 27804 49644 27860 49700
rect 27916 50764 27972 50820
rect 27804 48972 27860 49028
rect 28028 49756 28084 49812
rect 27356 48914 27412 48916
rect 27356 48862 27358 48914
rect 27358 48862 27410 48914
rect 27410 48862 27412 48914
rect 27356 48860 27412 48862
rect 27468 48300 27524 48356
rect 27244 48242 27300 48244
rect 27244 48190 27246 48242
rect 27246 48190 27298 48242
rect 27298 48190 27300 48242
rect 27244 48188 27300 48190
rect 27244 47570 27300 47572
rect 27244 47518 27246 47570
rect 27246 47518 27298 47570
rect 27298 47518 27300 47570
rect 27244 47516 27300 47518
rect 28028 48748 28084 48804
rect 27692 48188 27748 48244
rect 27468 46956 27524 47012
rect 27580 47964 27636 48020
rect 27468 46786 27524 46788
rect 27468 46734 27470 46786
rect 27470 46734 27522 46786
rect 27522 46734 27524 46786
rect 27468 46732 27524 46734
rect 27020 46396 27076 46452
rect 27468 46396 27524 46452
rect 27020 45778 27076 45780
rect 27020 45726 27022 45778
rect 27022 45726 27074 45778
rect 27074 45726 27076 45778
rect 27020 45724 27076 45726
rect 26908 45388 26964 45444
rect 27356 45612 27412 45668
rect 26796 44322 26852 44324
rect 26796 44270 26798 44322
rect 26798 44270 26850 44322
rect 26850 44270 26852 44322
rect 26796 44268 26852 44270
rect 26124 43596 26180 43652
rect 26348 43372 26404 43428
rect 25900 43148 25956 43204
rect 25564 42082 25620 42084
rect 25564 42030 25566 42082
rect 25566 42030 25618 42082
rect 25618 42030 25620 42082
rect 25564 42028 25620 42030
rect 25340 40796 25396 40852
rect 25676 41858 25732 41860
rect 25676 41806 25678 41858
rect 25678 41806 25730 41858
rect 25730 41806 25732 41858
rect 25676 41804 25732 41806
rect 25564 41020 25620 41076
rect 25676 40962 25732 40964
rect 25676 40910 25678 40962
rect 25678 40910 25730 40962
rect 25730 40910 25732 40962
rect 25676 40908 25732 40910
rect 26348 42812 26404 42868
rect 25900 42028 25956 42084
rect 26348 42252 26404 42308
rect 26012 41410 26068 41412
rect 26012 41358 26014 41410
rect 26014 41358 26066 41410
rect 26066 41358 26068 41410
rect 26012 41356 26068 41358
rect 26572 42866 26628 42868
rect 26572 42814 26574 42866
rect 26574 42814 26626 42866
rect 26626 42814 26628 42866
rect 26572 42812 26628 42814
rect 26796 43484 26852 43540
rect 27356 45388 27412 45444
rect 27020 44044 27076 44100
rect 27020 43650 27076 43652
rect 27020 43598 27022 43650
rect 27022 43598 27074 43650
rect 27074 43598 27076 43650
rect 27020 43596 27076 43598
rect 26908 42252 26964 42308
rect 26572 41692 26628 41748
rect 26796 42140 26852 42196
rect 27468 44828 27524 44884
rect 27692 47628 27748 47684
rect 27692 46844 27748 46900
rect 27692 45388 27748 45444
rect 28028 48300 28084 48356
rect 28028 47346 28084 47348
rect 28028 47294 28030 47346
rect 28030 47294 28082 47346
rect 28082 47294 28084 47346
rect 28028 47292 28084 47294
rect 27916 47068 27972 47124
rect 28028 45948 28084 46004
rect 28028 44994 28084 44996
rect 28028 44942 28030 44994
rect 28030 44942 28082 44994
rect 28082 44942 28084 44994
rect 28028 44940 28084 44942
rect 27804 44156 27860 44212
rect 27468 43036 27524 43092
rect 27580 43596 27636 43652
rect 27468 42866 27524 42868
rect 27468 42814 27470 42866
rect 27470 42814 27522 42866
rect 27522 42814 27524 42866
rect 27468 42812 27524 42814
rect 29260 55074 29316 55076
rect 29260 55022 29262 55074
rect 29262 55022 29314 55074
rect 29314 55022 29316 55074
rect 29260 55020 29316 55022
rect 29820 55020 29876 55076
rect 29596 53900 29652 53956
rect 28252 52556 28308 52612
rect 29148 53618 29204 53620
rect 29148 53566 29150 53618
rect 29150 53566 29202 53618
rect 29202 53566 29204 53618
rect 29148 53564 29204 53566
rect 29596 53564 29652 53620
rect 29036 53004 29092 53060
rect 28924 52834 28980 52836
rect 28924 52782 28926 52834
rect 28926 52782 28978 52834
rect 28978 52782 28980 52834
rect 28924 52780 28980 52782
rect 28588 52556 28644 52612
rect 28476 52444 28532 52500
rect 29484 53116 29540 53172
rect 30156 54348 30212 54404
rect 30380 54572 30436 54628
rect 30268 54236 30324 54292
rect 30380 54124 30436 54180
rect 29932 53900 29988 53956
rect 30156 53730 30212 53732
rect 30156 53678 30158 53730
rect 30158 53678 30210 53730
rect 30210 53678 30212 53730
rect 30156 53676 30212 53678
rect 29820 53340 29876 53396
rect 30716 56082 30772 56084
rect 30716 56030 30718 56082
rect 30718 56030 30770 56082
rect 30770 56030 30772 56082
rect 30716 56028 30772 56030
rect 36316 57708 36372 57764
rect 34300 56252 34356 56308
rect 30940 55916 30996 55972
rect 31052 55132 31108 55188
rect 32396 55970 32452 55972
rect 32396 55918 32398 55970
rect 32398 55918 32450 55970
rect 32450 55918 32452 55970
rect 32396 55916 32452 55918
rect 34300 55916 34356 55972
rect 31612 55468 31668 55524
rect 30604 54236 30660 54292
rect 31500 54402 31556 54404
rect 31500 54350 31502 54402
rect 31502 54350 31554 54402
rect 31554 54350 31556 54402
rect 31500 54348 31556 54350
rect 30940 53452 30996 53508
rect 31164 53788 31220 53844
rect 31164 53452 31220 53508
rect 31724 55356 31780 55412
rect 31724 55074 31780 55076
rect 31724 55022 31726 55074
rect 31726 55022 31778 55074
rect 31778 55022 31780 55074
rect 31724 55020 31780 55022
rect 31836 54290 31892 54292
rect 31836 54238 31838 54290
rect 31838 54238 31890 54290
rect 31890 54238 31892 54290
rect 31836 54236 31892 54238
rect 31724 53506 31780 53508
rect 31724 53454 31726 53506
rect 31726 53454 31778 53506
rect 31778 53454 31780 53506
rect 31724 53452 31780 53454
rect 31612 53340 31668 53396
rect 30604 53228 30660 53284
rect 31164 53116 31220 53172
rect 30716 53004 30772 53060
rect 29036 51660 29092 51716
rect 29372 50988 29428 51044
rect 28252 49756 28308 49812
rect 28252 49196 28308 49252
rect 28364 49420 28420 49476
rect 28924 49420 28980 49476
rect 29372 50316 29428 50372
rect 28364 49026 28420 49028
rect 28364 48974 28366 49026
rect 28366 48974 28418 49026
rect 28418 48974 28420 49026
rect 28364 48972 28420 48974
rect 28588 48972 28644 49028
rect 28476 48802 28532 48804
rect 28476 48750 28478 48802
rect 28478 48750 28530 48802
rect 28530 48750 28532 48802
rect 28476 48748 28532 48750
rect 29708 51938 29764 51940
rect 29708 51886 29710 51938
rect 29710 51886 29762 51938
rect 29762 51886 29764 51938
rect 29708 51884 29764 51886
rect 30380 51938 30436 51940
rect 30380 51886 30382 51938
rect 30382 51886 30434 51938
rect 30434 51886 30436 51938
rect 30380 51884 30436 51886
rect 29596 50092 29652 50148
rect 29372 49810 29428 49812
rect 29372 49758 29374 49810
rect 29374 49758 29426 49810
rect 29426 49758 29428 49810
rect 29372 49756 29428 49758
rect 29932 51548 29988 51604
rect 30156 51548 30212 51604
rect 29820 51100 29876 51156
rect 30044 50876 30100 50932
rect 30156 50818 30212 50820
rect 30156 50766 30158 50818
rect 30158 50766 30210 50818
rect 30210 50766 30212 50818
rect 30156 50764 30212 50766
rect 30044 50540 30100 50596
rect 30268 50540 30324 50596
rect 29484 49644 29540 49700
rect 29260 48972 29316 49028
rect 28252 48524 28308 48580
rect 28812 48748 28868 48804
rect 28588 48130 28644 48132
rect 28588 48078 28590 48130
rect 28590 48078 28642 48130
rect 28642 48078 28644 48130
rect 28588 48076 28644 48078
rect 29036 48748 29092 48804
rect 28364 47404 28420 47460
rect 28252 47068 28308 47124
rect 28252 45948 28308 46004
rect 28700 46956 28756 47012
rect 28588 46508 28644 46564
rect 28700 46620 28756 46676
rect 28588 46060 28644 46116
rect 28700 45724 28756 45780
rect 28924 46844 28980 46900
rect 28812 45500 28868 45556
rect 28924 45724 28980 45780
rect 28364 45164 28420 45220
rect 28476 45106 28532 45108
rect 28476 45054 28478 45106
rect 28478 45054 28530 45106
rect 28530 45054 28532 45106
rect 28476 45052 28532 45054
rect 28588 44492 28644 44548
rect 28812 45106 28868 45108
rect 28812 45054 28814 45106
rect 28814 45054 28866 45106
rect 28866 45054 28868 45106
rect 28812 45052 28868 45054
rect 29260 48636 29316 48692
rect 29820 48748 29876 48804
rect 29596 48412 29652 48468
rect 29820 48466 29876 48468
rect 29820 48414 29822 48466
rect 29822 48414 29874 48466
rect 29874 48414 29876 48466
rect 29820 48412 29876 48414
rect 29372 48188 29428 48244
rect 29596 47570 29652 47572
rect 29596 47518 29598 47570
rect 29598 47518 29650 47570
rect 29650 47518 29652 47570
rect 29596 47516 29652 47518
rect 29148 47068 29204 47124
rect 29260 46674 29316 46676
rect 29260 46622 29262 46674
rect 29262 46622 29314 46674
rect 29314 46622 29316 46674
rect 29260 46620 29316 46622
rect 29260 46284 29316 46340
rect 29036 44716 29092 44772
rect 29708 47346 29764 47348
rect 29708 47294 29710 47346
rect 29710 47294 29762 47346
rect 29762 47294 29764 47346
rect 29708 47292 29764 47294
rect 29820 46956 29876 47012
rect 29372 45948 29428 46004
rect 29596 46844 29652 46900
rect 29596 46396 29652 46452
rect 30380 49922 30436 49924
rect 30380 49870 30382 49922
rect 30382 49870 30434 49922
rect 30434 49870 30436 49922
rect 30380 49868 30436 49870
rect 30156 49420 30212 49476
rect 30268 48802 30324 48804
rect 30268 48750 30270 48802
rect 30270 48750 30322 48802
rect 30322 48750 30324 48802
rect 30268 48748 30324 48750
rect 30828 52162 30884 52164
rect 30828 52110 30830 52162
rect 30830 52110 30882 52162
rect 30882 52110 30884 52162
rect 30828 52108 30884 52110
rect 31948 53170 32004 53172
rect 31948 53118 31950 53170
rect 31950 53118 32002 53170
rect 32002 53118 32004 53170
rect 31948 53116 32004 53118
rect 31836 52668 31892 52724
rect 32732 55186 32788 55188
rect 32732 55134 32734 55186
rect 32734 55134 32786 55186
rect 32786 55134 32788 55186
rect 32732 55132 32788 55134
rect 32172 53618 32228 53620
rect 32172 53566 32174 53618
rect 32174 53566 32226 53618
rect 32226 53566 32228 53618
rect 32172 53564 32228 53566
rect 33180 55132 33236 55188
rect 33180 53900 33236 53956
rect 32956 53676 33012 53732
rect 32060 52556 32116 52612
rect 33292 53564 33348 53620
rect 31836 52274 31892 52276
rect 31836 52222 31838 52274
rect 31838 52222 31890 52274
rect 31890 52222 31892 52274
rect 31836 52220 31892 52222
rect 30604 51548 30660 51604
rect 30716 50764 30772 50820
rect 33068 52668 33124 52724
rect 31276 51378 31332 51380
rect 31276 51326 31278 51378
rect 31278 51326 31330 51378
rect 31330 51326 31332 51378
rect 31276 51324 31332 51326
rect 31164 50764 31220 50820
rect 31612 50988 31668 51044
rect 30604 50428 30660 50484
rect 31052 50594 31108 50596
rect 31052 50542 31054 50594
rect 31054 50542 31106 50594
rect 31106 50542 31108 50594
rect 31052 50540 31108 50542
rect 31388 50482 31444 50484
rect 31388 50430 31390 50482
rect 31390 50430 31442 50482
rect 31442 50430 31444 50482
rect 31388 50428 31444 50430
rect 32060 51154 32116 51156
rect 32060 51102 32062 51154
rect 32062 51102 32114 51154
rect 32114 51102 32116 51154
rect 32060 51100 32116 51102
rect 32284 50988 32340 51044
rect 32284 50652 32340 50708
rect 32172 50428 32228 50484
rect 32956 51548 33012 51604
rect 30716 50204 30772 50260
rect 31724 50092 31780 50148
rect 31276 49922 31332 49924
rect 31276 49870 31278 49922
rect 31278 49870 31330 49922
rect 31330 49870 31332 49922
rect 31276 49868 31332 49870
rect 30828 49756 30884 49812
rect 31388 49756 31444 49812
rect 30828 49084 30884 49140
rect 30940 49420 30996 49476
rect 30716 48972 30772 49028
rect 30268 48412 30324 48468
rect 30268 48242 30324 48244
rect 30268 48190 30270 48242
rect 30270 48190 30322 48242
rect 30322 48190 30324 48242
rect 30268 48188 30324 48190
rect 30156 47068 30212 47124
rect 30044 46844 30100 46900
rect 30156 46786 30212 46788
rect 30156 46734 30158 46786
rect 30158 46734 30210 46786
rect 30210 46734 30212 46786
rect 30156 46732 30212 46734
rect 30492 47682 30548 47684
rect 30492 47630 30494 47682
rect 30494 47630 30546 47682
rect 30546 47630 30548 47682
rect 30492 47628 30548 47630
rect 30380 47346 30436 47348
rect 30380 47294 30382 47346
rect 30382 47294 30434 47346
rect 30434 47294 30436 47346
rect 30380 47292 30436 47294
rect 29932 46284 29988 46340
rect 30268 46284 30324 46340
rect 30044 46002 30100 46004
rect 30044 45950 30046 46002
rect 30046 45950 30098 46002
rect 30098 45950 30100 46002
rect 30044 45948 30100 45950
rect 29484 45836 29540 45892
rect 29260 45500 29316 45556
rect 29932 45388 29988 45444
rect 29708 45218 29764 45220
rect 29708 45166 29710 45218
rect 29710 45166 29762 45218
rect 29762 45166 29764 45218
rect 29708 45164 29764 45166
rect 28700 44380 28756 44436
rect 29260 44546 29316 44548
rect 29260 44494 29262 44546
rect 29262 44494 29314 44546
rect 29314 44494 29316 44546
rect 29260 44492 29316 44494
rect 29372 44380 29428 44436
rect 29484 44322 29540 44324
rect 29484 44270 29486 44322
rect 29486 44270 29538 44322
rect 29538 44270 29540 44322
rect 29484 44268 29540 44270
rect 27580 42754 27636 42756
rect 27580 42702 27582 42754
rect 27582 42702 27634 42754
rect 27634 42702 27636 42754
rect 27580 42700 27636 42702
rect 26460 41580 26516 41636
rect 26348 41356 26404 41412
rect 26124 40962 26180 40964
rect 26124 40910 26126 40962
rect 26126 40910 26178 40962
rect 26178 40910 26180 40962
rect 26124 40908 26180 40910
rect 25452 39564 25508 39620
rect 25564 40236 25620 40292
rect 25340 39452 25396 39508
rect 24892 38556 24948 38612
rect 24220 37772 24276 37828
rect 23996 37490 24052 37492
rect 23996 37438 23998 37490
rect 23998 37438 24050 37490
rect 24050 37438 24052 37490
rect 23996 37436 24052 37438
rect 24332 37490 24388 37492
rect 24332 37438 24334 37490
rect 24334 37438 24386 37490
rect 24386 37438 24388 37490
rect 24332 37436 24388 37438
rect 25340 37324 25396 37380
rect 23996 36316 24052 36372
rect 23660 34300 23716 34356
rect 24332 35868 24388 35924
rect 24668 35980 24724 36036
rect 24220 33964 24276 34020
rect 24780 34914 24836 34916
rect 24780 34862 24782 34914
rect 24782 34862 24834 34914
rect 24834 34862 24836 34914
rect 24780 34860 24836 34862
rect 23436 33516 23492 33572
rect 25788 40402 25844 40404
rect 25788 40350 25790 40402
rect 25790 40350 25842 40402
rect 25842 40350 25844 40402
rect 25788 40348 25844 40350
rect 26012 39788 26068 39844
rect 25676 39004 25732 39060
rect 26012 39004 26068 39060
rect 25340 35980 25396 36036
rect 26124 38780 26180 38836
rect 25676 36258 25732 36260
rect 25676 36206 25678 36258
rect 25678 36206 25730 36258
rect 25730 36206 25732 36258
rect 25676 36204 25732 36206
rect 26012 37826 26068 37828
rect 26012 37774 26014 37826
rect 26014 37774 26066 37826
rect 26066 37774 26068 37826
rect 26012 37772 26068 37774
rect 26236 38220 26292 38276
rect 26236 37548 26292 37604
rect 27356 41970 27412 41972
rect 27356 41918 27358 41970
rect 27358 41918 27410 41970
rect 27410 41918 27412 41970
rect 27356 41916 27412 41918
rect 27020 41804 27076 41860
rect 26572 40626 26628 40628
rect 26572 40574 26574 40626
rect 26574 40574 26626 40626
rect 26626 40574 26628 40626
rect 26572 40572 26628 40574
rect 27132 40514 27188 40516
rect 27132 40462 27134 40514
rect 27134 40462 27186 40514
rect 27186 40462 27188 40514
rect 27132 40460 27188 40462
rect 27244 40236 27300 40292
rect 26796 39004 26852 39060
rect 26908 39340 26964 39396
rect 27804 43036 27860 43092
rect 27916 42364 27972 42420
rect 27804 41356 27860 41412
rect 27692 40236 27748 40292
rect 27580 39788 27636 39844
rect 27692 39676 27748 39732
rect 27468 38780 27524 38836
rect 26572 38050 26628 38052
rect 26572 37998 26574 38050
rect 26574 37998 26626 38050
rect 26626 37998 26628 38050
rect 26572 37996 26628 37998
rect 26572 37548 26628 37604
rect 26908 37826 26964 37828
rect 26908 37774 26910 37826
rect 26910 37774 26962 37826
rect 26962 37774 26964 37826
rect 26908 37772 26964 37774
rect 26796 37660 26852 37716
rect 26908 37324 26964 37380
rect 27132 37884 27188 37940
rect 26236 36706 26292 36708
rect 26236 36654 26238 36706
rect 26238 36654 26290 36706
rect 26290 36654 26292 36706
rect 26236 36652 26292 36654
rect 26572 36594 26628 36596
rect 26572 36542 26574 36594
rect 26574 36542 26626 36594
rect 26626 36542 26628 36594
rect 26572 36540 26628 36542
rect 26460 36428 26516 36484
rect 26684 36204 26740 36260
rect 27916 40572 27972 40628
rect 28252 42476 28308 42532
rect 28588 43596 28644 43652
rect 29148 43650 29204 43652
rect 29148 43598 29150 43650
rect 29150 43598 29202 43650
rect 29202 43598 29204 43650
rect 29148 43596 29204 43598
rect 28588 43314 28644 43316
rect 28588 43262 28590 43314
rect 28590 43262 28642 43314
rect 28642 43262 28644 43314
rect 28588 43260 28644 43262
rect 28924 43148 28980 43204
rect 28364 41916 28420 41972
rect 28700 42754 28756 42756
rect 28700 42702 28702 42754
rect 28702 42702 28754 42754
rect 28754 42702 28756 42754
rect 28700 42700 28756 42702
rect 29036 43036 29092 43092
rect 28924 42082 28980 42084
rect 28924 42030 28926 42082
rect 28926 42030 28978 42082
rect 28978 42030 28980 42082
rect 28924 42028 28980 42030
rect 28476 41692 28532 41748
rect 28028 39730 28084 39732
rect 28028 39678 28030 39730
rect 28030 39678 28082 39730
rect 28082 39678 28084 39730
rect 28028 39676 28084 39678
rect 28028 39340 28084 39396
rect 28364 40572 28420 40628
rect 28700 41074 28756 41076
rect 28700 41022 28702 41074
rect 28702 41022 28754 41074
rect 28754 41022 28756 41074
rect 28700 41020 28756 41022
rect 29036 40908 29092 40964
rect 28588 40514 28644 40516
rect 28588 40462 28590 40514
rect 28590 40462 28642 40514
rect 28642 40462 28644 40514
rect 28588 40460 28644 40462
rect 28588 39394 28644 39396
rect 28588 39342 28590 39394
rect 28590 39342 28642 39394
rect 28642 39342 28644 39394
rect 28588 39340 28644 39342
rect 27692 37660 27748 37716
rect 27804 37436 27860 37492
rect 27468 36988 27524 37044
rect 27804 36988 27860 37044
rect 28140 38108 28196 38164
rect 28252 37884 28308 37940
rect 28028 37772 28084 37828
rect 27356 36316 27412 36372
rect 26684 35980 26740 36036
rect 27356 35980 27412 36036
rect 27356 35644 27412 35700
rect 26348 35308 26404 35364
rect 25900 35026 25956 35028
rect 25900 34974 25902 35026
rect 25902 34974 25954 35026
rect 25954 34974 25956 35026
rect 25900 34972 25956 34974
rect 26684 34972 26740 35028
rect 26348 34914 26404 34916
rect 26348 34862 26350 34914
rect 26350 34862 26402 34914
rect 26402 34862 26404 34914
rect 26348 34860 26404 34862
rect 25564 34748 25620 34804
rect 27244 34914 27300 34916
rect 27244 34862 27246 34914
rect 27246 34862 27298 34914
rect 27298 34862 27300 34914
rect 27244 34860 27300 34862
rect 27580 36482 27636 36484
rect 27580 36430 27582 36482
rect 27582 36430 27634 36482
rect 27634 36430 27636 36482
rect 27580 36428 27636 36430
rect 24892 34412 24948 34468
rect 25676 34242 25732 34244
rect 25676 34190 25678 34242
rect 25678 34190 25730 34242
rect 25730 34190 25732 34242
rect 25676 34188 25732 34190
rect 25564 34130 25620 34132
rect 25564 34078 25566 34130
rect 25566 34078 25618 34130
rect 25618 34078 25620 34130
rect 25564 34076 25620 34078
rect 25676 33852 25732 33908
rect 26236 34354 26292 34356
rect 26236 34302 26238 34354
rect 26238 34302 26290 34354
rect 26290 34302 26292 34354
rect 26236 34300 26292 34302
rect 26012 33852 26068 33908
rect 25004 33516 25060 33572
rect 21980 33346 22036 33348
rect 21980 33294 21982 33346
rect 21982 33294 22034 33346
rect 22034 33294 22036 33346
rect 21980 33292 22036 33294
rect 22092 33234 22148 33236
rect 22092 33182 22094 33234
rect 22094 33182 22146 33234
rect 22146 33182 22148 33234
rect 22092 33180 22148 33182
rect 24332 33404 24388 33460
rect 23996 33122 24052 33124
rect 23996 33070 23998 33122
rect 23998 33070 24050 33122
rect 24050 33070 24052 33122
rect 23996 33068 24052 33070
rect 25676 33346 25732 33348
rect 25676 33294 25678 33346
rect 25678 33294 25730 33346
rect 25730 33294 25732 33346
rect 25676 33292 25732 33294
rect 24444 33180 24500 33236
rect 25564 33180 25620 33236
rect 24780 33068 24836 33124
rect 25452 33068 25508 33124
rect 23436 32674 23492 32676
rect 23436 32622 23438 32674
rect 23438 32622 23490 32674
rect 23490 32622 23492 32674
rect 23436 32620 23492 32622
rect 25228 32674 25284 32676
rect 25228 32622 25230 32674
rect 25230 32622 25282 32674
rect 25282 32622 25284 32674
rect 25228 32620 25284 32622
rect 26348 34130 26404 34132
rect 26348 34078 26350 34130
rect 26350 34078 26402 34130
rect 26402 34078 26404 34130
rect 26348 34076 26404 34078
rect 25900 33068 25956 33124
rect 23100 32284 23156 32340
rect 23548 32338 23604 32340
rect 23548 32286 23550 32338
rect 23550 32286 23602 32338
rect 23602 32286 23604 32338
rect 23548 32284 23604 32286
rect 24220 32284 24276 32340
rect 21196 31836 21252 31892
rect 21980 31724 22036 31780
rect 21868 31106 21924 31108
rect 21868 31054 21870 31106
rect 21870 31054 21922 31106
rect 21922 31054 21924 31106
rect 21868 31052 21924 31054
rect 21308 30716 21364 30772
rect 21756 30828 21812 30884
rect 23996 30716 24052 30772
rect 21308 30098 21364 30100
rect 21308 30046 21310 30098
rect 21310 30046 21362 30098
rect 21362 30046 21364 30098
rect 21308 30044 21364 30046
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20636 29820 20692 29876
rect 20044 29764 20100 29766
rect 19964 29650 20020 29652
rect 19964 29598 19966 29650
rect 19966 29598 20018 29650
rect 20018 29598 20020 29650
rect 19964 29596 20020 29598
rect 20636 29596 20692 29652
rect 19852 29538 19908 29540
rect 19852 29486 19854 29538
rect 19854 29486 19906 29538
rect 19906 29486 19908 29538
rect 19852 29484 19908 29486
rect 17612 28588 17668 28644
rect 18508 29148 18564 29204
rect 18620 28924 18676 28980
rect 18956 29314 19012 29316
rect 18956 29262 18958 29314
rect 18958 29262 19010 29314
rect 19010 29262 19012 29314
rect 18956 29260 19012 29262
rect 19740 29314 19796 29316
rect 19740 29262 19742 29314
rect 19742 29262 19794 29314
rect 19794 29262 19796 29314
rect 19740 29260 19796 29262
rect 19292 28812 19348 28868
rect 17612 27916 17668 27972
rect 17388 27858 17444 27860
rect 17388 27806 17390 27858
rect 17390 27806 17442 27858
rect 17442 27806 17444 27858
rect 17388 27804 17444 27806
rect 17948 27746 18004 27748
rect 17948 27694 17950 27746
rect 17950 27694 18002 27746
rect 18002 27694 18004 27746
rect 17948 27692 18004 27694
rect 17612 27132 17668 27188
rect 17388 26236 17444 26292
rect 17836 26796 17892 26852
rect 17388 26012 17444 26068
rect 17500 25900 17556 25956
rect 16492 23100 16548 23156
rect 15820 22428 15876 22484
rect 15708 22146 15764 22148
rect 15708 22094 15710 22146
rect 15710 22094 15762 22146
rect 15762 22094 15764 22146
rect 15708 22092 15764 22094
rect 15148 20972 15204 21028
rect 15148 20130 15204 20132
rect 15148 20078 15150 20130
rect 15150 20078 15202 20130
rect 15202 20078 15204 20130
rect 15148 20076 15204 20078
rect 15036 19346 15092 19348
rect 15036 19294 15038 19346
rect 15038 19294 15090 19346
rect 15090 19294 15092 19346
rect 15036 19292 15092 19294
rect 14812 19180 14868 19236
rect 15036 19068 15092 19124
rect 14476 17442 14532 17444
rect 14476 17390 14478 17442
rect 14478 17390 14530 17442
rect 14530 17390 14532 17442
rect 14476 17388 14532 17390
rect 14476 17164 14532 17220
rect 14476 15932 14532 15988
rect 14588 16380 14644 16436
rect 14252 15484 14308 15540
rect 14252 15260 14308 15316
rect 14028 12962 14084 12964
rect 14028 12910 14030 12962
rect 14030 12910 14082 12962
rect 14082 12910 14084 12962
rect 14028 12908 14084 12910
rect 14028 12012 14084 12068
rect 13468 10444 13524 10500
rect 13580 10556 13636 10612
rect 13804 9772 13860 9828
rect 13692 9660 13748 9716
rect 14028 11004 14084 11060
rect 14588 14588 14644 14644
rect 14476 14140 14532 14196
rect 14924 16940 14980 16996
rect 14924 16492 14980 16548
rect 15372 20748 15428 20804
rect 15260 18172 15316 18228
rect 15820 20076 15876 20132
rect 15596 19852 15652 19908
rect 15708 19122 15764 19124
rect 15708 19070 15710 19122
rect 15710 19070 15762 19122
rect 15762 19070 15764 19122
rect 15708 19068 15764 19070
rect 15148 17052 15204 17108
rect 15820 17778 15876 17780
rect 15820 17726 15822 17778
rect 15822 17726 15874 17778
rect 15874 17726 15876 17778
rect 15820 17724 15876 17726
rect 15932 17836 15988 17892
rect 15484 17500 15540 17556
rect 15372 17052 15428 17108
rect 15372 16828 15428 16884
rect 15036 16380 15092 16436
rect 14924 16268 14980 16324
rect 15260 16210 15316 16212
rect 15260 16158 15262 16210
rect 15262 16158 15314 16210
rect 15314 16158 15316 16210
rect 15260 16156 15316 16158
rect 14924 15372 14980 15428
rect 14924 14140 14980 14196
rect 15260 15090 15316 15092
rect 15260 15038 15262 15090
rect 15262 15038 15314 15090
rect 15314 15038 15316 15090
rect 15260 15036 15316 15038
rect 15484 16156 15540 16212
rect 15932 17164 15988 17220
rect 16828 23826 16884 23828
rect 16828 23774 16830 23826
rect 16830 23774 16882 23826
rect 16882 23774 16884 23826
rect 16828 23772 16884 23774
rect 16940 23660 16996 23716
rect 16940 23436 16996 23492
rect 16716 23100 16772 23156
rect 17836 25564 17892 25620
rect 17500 25452 17556 25508
rect 18060 27074 18116 27076
rect 18060 27022 18062 27074
rect 18062 27022 18114 27074
rect 18114 27022 18116 27074
rect 18060 27020 18116 27022
rect 19740 28642 19796 28644
rect 19740 28590 19742 28642
rect 19742 28590 19794 28642
rect 19794 28590 19796 28642
rect 19740 28588 19796 28590
rect 20524 28588 20580 28644
rect 18956 28476 19012 28532
rect 20300 28418 20356 28420
rect 20300 28366 20302 28418
rect 20302 28366 20354 28418
rect 20354 28366 20356 28418
rect 20300 28364 20356 28366
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 18060 26124 18116 26180
rect 18172 26236 18228 26292
rect 19404 27692 19460 27748
rect 18732 26572 18788 26628
rect 18620 26290 18676 26292
rect 18620 26238 18622 26290
rect 18622 26238 18674 26290
rect 18674 26238 18676 26290
rect 18620 26236 18676 26238
rect 18284 26124 18340 26180
rect 18172 25564 18228 25620
rect 17388 24108 17444 24164
rect 17388 23772 17444 23828
rect 17052 22988 17108 23044
rect 17276 23324 17332 23380
rect 17724 25394 17780 25396
rect 17724 25342 17726 25394
rect 17726 25342 17778 25394
rect 17778 25342 17780 25394
rect 17724 25340 17780 25342
rect 17836 25228 17892 25284
rect 17612 24220 17668 24276
rect 17724 24668 17780 24724
rect 17836 24108 17892 24164
rect 18172 23996 18228 24052
rect 17612 23378 17668 23380
rect 17612 23326 17614 23378
rect 17614 23326 17666 23378
rect 17666 23326 17668 23378
rect 17612 23324 17668 23326
rect 18060 23154 18116 23156
rect 18060 23102 18062 23154
rect 18062 23102 18114 23154
rect 18114 23102 18116 23154
rect 18060 23100 18116 23102
rect 17276 22876 17332 22932
rect 17052 22652 17108 22708
rect 16716 22482 16772 22484
rect 16716 22430 16718 22482
rect 16718 22430 16770 22482
rect 16770 22430 16772 22482
rect 16716 22428 16772 22430
rect 16604 21868 16660 21924
rect 16156 21586 16212 21588
rect 16156 21534 16158 21586
rect 16158 21534 16210 21586
rect 16210 21534 16212 21586
rect 16156 21532 16212 21534
rect 16268 20300 16324 20356
rect 16716 20972 16772 21028
rect 18172 22764 18228 22820
rect 17724 21810 17780 21812
rect 17724 21758 17726 21810
rect 17726 21758 17778 21810
rect 17778 21758 17780 21810
rect 17724 21756 17780 21758
rect 18396 24220 18452 24276
rect 18508 24050 18564 24052
rect 18508 23998 18510 24050
rect 18510 23998 18562 24050
rect 18562 23998 18564 24050
rect 18508 23996 18564 23998
rect 18284 21474 18340 21476
rect 18284 21422 18286 21474
rect 18286 21422 18338 21474
rect 18338 21422 18340 21474
rect 18284 21420 18340 21422
rect 18172 21084 18228 21140
rect 16268 18562 16324 18564
rect 16268 18510 16270 18562
rect 16270 18510 16322 18562
rect 16322 18510 16324 18562
rect 16268 18508 16324 18510
rect 16156 17052 16212 17108
rect 15932 16828 15988 16884
rect 15484 15314 15540 15316
rect 15484 15262 15486 15314
rect 15486 15262 15538 15314
rect 15538 15262 15540 15314
rect 15484 15260 15540 15262
rect 15260 14530 15316 14532
rect 15260 14478 15262 14530
rect 15262 14478 15314 14530
rect 15314 14478 15316 14530
rect 15260 14476 15316 14478
rect 15484 14924 15540 14980
rect 14588 12796 14644 12852
rect 14252 9772 14308 9828
rect 13468 9212 13524 9268
rect 12236 6972 12292 7028
rect 11900 6636 11956 6692
rect 11900 5516 11956 5572
rect 12348 6130 12404 6132
rect 12348 6078 12350 6130
rect 12350 6078 12402 6130
rect 12402 6078 12404 6130
rect 12348 6076 12404 6078
rect 12684 6412 12740 6468
rect 12572 5516 12628 5572
rect 12796 5292 12852 5348
rect 13132 5628 13188 5684
rect 12012 3836 12068 3892
rect 11900 2828 11956 2884
rect 13916 9100 13972 9156
rect 13468 8428 13524 8484
rect 14028 8316 14084 8372
rect 13804 8258 13860 8260
rect 13804 8206 13806 8258
rect 13806 8206 13858 8258
rect 13858 8206 13860 8258
rect 13804 8204 13860 8206
rect 13356 8092 13412 8148
rect 13468 7474 13524 7476
rect 13468 7422 13470 7474
rect 13470 7422 13522 7474
rect 13522 7422 13524 7474
rect 13468 7420 13524 7422
rect 13580 7308 13636 7364
rect 14028 6914 14084 6916
rect 14028 6862 14030 6914
rect 14030 6862 14082 6914
rect 14082 6862 14084 6914
rect 14028 6860 14084 6862
rect 14476 9324 14532 9380
rect 14364 9266 14420 9268
rect 14364 9214 14366 9266
rect 14366 9214 14418 9266
rect 14418 9214 14420 9266
rect 14364 9212 14420 9214
rect 14364 8258 14420 8260
rect 14364 8206 14366 8258
rect 14366 8206 14418 8258
rect 14418 8206 14420 8258
rect 14364 8204 14420 8206
rect 14700 9938 14756 9940
rect 14700 9886 14702 9938
rect 14702 9886 14754 9938
rect 14754 9886 14756 9938
rect 14700 9884 14756 9886
rect 14924 13746 14980 13748
rect 14924 13694 14926 13746
rect 14926 13694 14978 13746
rect 14978 13694 14980 13746
rect 14924 13692 14980 13694
rect 15036 13132 15092 13188
rect 15148 13186 15204 13188
rect 15148 13134 15150 13186
rect 15150 13134 15202 13186
rect 15202 13134 15204 13186
rect 15148 13132 15204 13134
rect 15372 12460 15428 12516
rect 15260 12348 15316 12404
rect 15596 13132 15652 13188
rect 15484 11788 15540 11844
rect 15372 10332 15428 10388
rect 14588 7586 14644 7588
rect 14588 7534 14590 7586
rect 14590 7534 14642 7586
rect 14642 7534 14644 7586
rect 14588 7532 14644 7534
rect 14924 9996 14980 10052
rect 13468 6748 13524 6804
rect 13468 5516 13524 5572
rect 13692 6636 13748 6692
rect 14812 9324 14868 9380
rect 14924 9154 14980 9156
rect 14924 9102 14926 9154
rect 14926 9102 14978 9154
rect 14978 9102 14980 9154
rect 14924 9100 14980 9102
rect 15708 11564 15764 11620
rect 15596 10668 15652 10724
rect 15372 8204 15428 8260
rect 15484 9212 15540 9268
rect 15260 7868 15316 7924
rect 15372 7980 15428 8036
rect 15932 14364 15988 14420
rect 15932 12572 15988 12628
rect 15708 10332 15764 10388
rect 15820 11228 15876 11284
rect 16604 20636 16660 20692
rect 16716 20524 16772 20580
rect 16716 19964 16772 20020
rect 16604 19628 16660 19684
rect 16604 19404 16660 19460
rect 16604 18956 16660 19012
rect 17612 20802 17668 20804
rect 17612 20750 17614 20802
rect 17614 20750 17666 20802
rect 17666 20750 17668 20802
rect 17612 20748 17668 20750
rect 17724 20412 17780 20468
rect 17948 20748 18004 20804
rect 17388 20300 17444 20356
rect 17836 20300 17892 20356
rect 16940 19964 16996 20020
rect 17612 19964 17668 20020
rect 17500 19740 17556 19796
rect 17164 19404 17220 19460
rect 17164 19068 17220 19124
rect 16828 18620 16884 18676
rect 16716 18562 16772 18564
rect 16716 18510 16718 18562
rect 16718 18510 16770 18562
rect 16770 18510 16772 18562
rect 16716 18508 16772 18510
rect 16604 18060 16660 18116
rect 17500 19068 17556 19124
rect 17276 18284 17332 18340
rect 16940 18060 16996 18116
rect 16940 17612 16996 17668
rect 18060 20130 18116 20132
rect 18060 20078 18062 20130
rect 18062 20078 18114 20130
rect 18114 20078 18116 20130
rect 18060 20076 18116 20078
rect 17612 18396 17668 18452
rect 17276 17500 17332 17556
rect 16604 17276 16660 17332
rect 16492 16210 16548 16212
rect 16492 16158 16494 16210
rect 16494 16158 16546 16210
rect 16546 16158 16548 16210
rect 16492 16156 16548 16158
rect 16828 16882 16884 16884
rect 16828 16830 16830 16882
rect 16830 16830 16882 16882
rect 16882 16830 16884 16882
rect 16828 16828 16884 16830
rect 16828 16492 16884 16548
rect 17724 18338 17780 18340
rect 17724 18286 17726 18338
rect 17726 18286 17778 18338
rect 17778 18286 17780 18338
rect 17724 18284 17780 18286
rect 17612 17948 17668 18004
rect 17388 17276 17444 17332
rect 17724 17666 17780 17668
rect 17724 17614 17726 17666
rect 17726 17614 17778 17666
rect 17778 17614 17780 17666
rect 17724 17612 17780 17614
rect 17612 17164 17668 17220
rect 17724 17388 17780 17444
rect 17500 16380 17556 16436
rect 16940 16044 16996 16100
rect 16940 15820 16996 15876
rect 16268 13746 16324 13748
rect 16268 13694 16270 13746
rect 16270 13694 16322 13746
rect 16322 13694 16324 13746
rect 16268 13692 16324 13694
rect 16604 12684 16660 12740
rect 16380 12460 16436 12516
rect 16156 11676 16212 11732
rect 16156 10556 16212 10612
rect 15932 9548 15988 9604
rect 15596 8652 15652 8708
rect 15708 9324 15764 9380
rect 15820 9266 15876 9268
rect 15820 9214 15822 9266
rect 15822 9214 15874 9266
rect 15874 9214 15876 9266
rect 15820 9212 15876 9214
rect 15932 9100 15988 9156
rect 16716 11900 16772 11956
rect 16940 15372 16996 15428
rect 16716 11676 16772 11732
rect 16716 11228 16772 11284
rect 16156 8988 16212 9044
rect 15708 8540 15764 8596
rect 15820 8764 15876 8820
rect 15484 7644 15540 7700
rect 15484 7474 15540 7476
rect 15484 7422 15486 7474
rect 15486 7422 15538 7474
rect 15538 7422 15540 7474
rect 15484 7420 15540 7422
rect 14476 6802 14532 6804
rect 14476 6750 14478 6802
rect 14478 6750 14530 6802
rect 14530 6750 14532 6802
rect 14476 6748 14532 6750
rect 14476 6076 14532 6132
rect 14700 6524 14756 6580
rect 14588 5682 14644 5684
rect 14588 5630 14590 5682
rect 14590 5630 14642 5682
rect 14642 5630 14644 5682
rect 14588 5628 14644 5630
rect 14028 5234 14084 5236
rect 14028 5182 14030 5234
rect 14030 5182 14082 5234
rect 14082 5182 14084 5234
rect 14028 5180 14084 5182
rect 14812 5346 14868 5348
rect 14812 5294 14814 5346
rect 14814 5294 14866 5346
rect 14866 5294 14868 5346
rect 14812 5292 14868 5294
rect 15148 5964 15204 6020
rect 16492 8540 16548 8596
rect 15932 8316 15988 8372
rect 16380 8316 16436 8372
rect 16268 8258 16324 8260
rect 16268 8206 16270 8258
rect 16270 8206 16322 8258
rect 16322 8206 16324 8258
rect 16268 8204 16324 8206
rect 16156 8092 16212 8148
rect 15932 7644 15988 7700
rect 15708 6524 15764 6580
rect 15596 5852 15652 5908
rect 14364 4956 14420 5012
rect 14700 3836 14756 3892
rect 15260 5068 15316 5124
rect 15820 6412 15876 6468
rect 16156 7420 16212 7476
rect 16268 7362 16324 7364
rect 16268 7310 16270 7362
rect 16270 7310 16322 7362
rect 16322 7310 16324 7362
rect 16268 7308 16324 7310
rect 16940 13580 16996 13636
rect 17164 16210 17220 16212
rect 17164 16158 17166 16210
rect 17166 16158 17218 16210
rect 17218 16158 17220 16210
rect 17164 16156 17220 16158
rect 17948 17276 18004 17332
rect 17948 17052 18004 17108
rect 17948 16828 18004 16884
rect 18620 21980 18676 22036
rect 18620 21586 18676 21588
rect 18620 21534 18622 21586
rect 18622 21534 18674 21586
rect 18674 21534 18676 21586
rect 18620 21532 18676 21534
rect 19404 26684 19460 26740
rect 19852 27356 19908 27412
rect 19628 26684 19684 26740
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19852 26348 19908 26404
rect 18844 26236 18900 26292
rect 19740 26236 19796 26292
rect 19068 26124 19124 26180
rect 18956 24444 19012 24500
rect 19516 25564 19572 25620
rect 20188 26290 20244 26292
rect 20188 26238 20190 26290
rect 20190 26238 20242 26290
rect 20242 26238 20244 26290
rect 20188 26236 20244 26238
rect 21196 29596 21252 29652
rect 20748 29314 20804 29316
rect 20748 29262 20750 29314
rect 20750 29262 20802 29314
rect 20802 29262 20804 29314
rect 20748 29260 20804 29262
rect 21308 29260 21364 29316
rect 21756 29986 21812 29988
rect 21756 29934 21758 29986
rect 21758 29934 21810 29986
rect 21810 29934 21812 29986
rect 21756 29932 21812 29934
rect 21980 29650 22036 29652
rect 21980 29598 21982 29650
rect 21982 29598 22034 29650
rect 22034 29598 22036 29650
rect 21980 29596 22036 29598
rect 21644 29260 21700 29316
rect 22316 30156 22372 30212
rect 22204 29538 22260 29540
rect 22204 29486 22206 29538
rect 22206 29486 22258 29538
rect 22258 29486 22260 29538
rect 22204 29484 22260 29486
rect 23772 30210 23828 30212
rect 23772 30158 23774 30210
rect 23774 30158 23826 30210
rect 23826 30158 23828 30210
rect 23772 30156 23828 30158
rect 22540 29986 22596 29988
rect 22540 29934 22542 29986
rect 22542 29934 22594 29986
rect 22594 29934 22596 29986
rect 22540 29932 22596 29934
rect 21980 28700 22036 28756
rect 21644 28588 21700 28644
rect 20524 26402 20580 26404
rect 20524 26350 20526 26402
rect 20526 26350 20578 26402
rect 20578 26350 20580 26402
rect 20524 26348 20580 26350
rect 20412 26124 20468 26180
rect 19852 25676 19908 25732
rect 20188 25506 20244 25508
rect 20188 25454 20190 25506
rect 20190 25454 20242 25506
rect 20242 25454 20244 25506
rect 20188 25452 20244 25454
rect 19404 24780 19460 24836
rect 19404 23772 19460 23828
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20188 24722 20244 24724
rect 20188 24670 20190 24722
rect 20190 24670 20242 24722
rect 20242 24670 20244 24722
rect 20188 24668 20244 24670
rect 19292 22764 19348 22820
rect 19628 24108 19684 24164
rect 19180 22370 19236 22372
rect 19180 22318 19182 22370
rect 19182 22318 19234 22370
rect 19234 22318 19236 22370
rect 19180 22316 19236 22318
rect 18956 22204 19012 22260
rect 18844 21532 18900 21588
rect 18844 21308 18900 21364
rect 19068 21420 19124 21476
rect 18732 20748 18788 20804
rect 18956 21196 19012 21252
rect 18620 20018 18676 20020
rect 18620 19966 18622 20018
rect 18622 19966 18674 20018
rect 18674 19966 18676 20018
rect 18620 19964 18676 19966
rect 18396 19404 18452 19460
rect 18172 16940 18228 16996
rect 17948 16492 18004 16548
rect 17052 12348 17108 12404
rect 17164 11788 17220 11844
rect 16940 11452 16996 11508
rect 16940 11004 16996 11060
rect 16828 10780 16884 10836
rect 16940 10668 16996 10724
rect 17164 11228 17220 11284
rect 16716 9436 16772 9492
rect 17052 9772 17108 9828
rect 16940 9212 16996 9268
rect 17500 14588 17556 14644
rect 18060 16156 18116 16212
rect 17948 15260 18004 15316
rect 18172 15484 18228 15540
rect 18844 20412 18900 20468
rect 18620 18956 18676 19012
rect 18732 19234 18788 19236
rect 18732 19182 18734 19234
rect 18734 19182 18786 19234
rect 18786 19182 18788 19234
rect 18732 19180 18788 19182
rect 18620 18396 18676 18452
rect 18844 18508 18900 18564
rect 18732 17836 18788 17892
rect 18620 17388 18676 17444
rect 18508 17164 18564 17220
rect 20748 26850 20804 26852
rect 20748 26798 20750 26850
rect 20750 26798 20802 26850
rect 20802 26798 20804 26850
rect 20748 26796 20804 26798
rect 21532 28418 21588 28420
rect 21532 28366 21534 28418
rect 21534 28366 21586 28418
rect 21586 28366 21588 28418
rect 21532 28364 21588 28366
rect 21532 27356 21588 27412
rect 21308 26962 21364 26964
rect 21308 26910 21310 26962
rect 21310 26910 21362 26962
rect 21362 26910 21364 26962
rect 21308 26908 21364 26910
rect 20860 26348 20916 26404
rect 20860 25676 20916 25732
rect 22316 28364 22372 28420
rect 22316 27916 22372 27972
rect 23996 29596 24052 29652
rect 22876 29314 22932 29316
rect 22876 29262 22878 29314
rect 22878 29262 22930 29314
rect 22930 29262 22932 29314
rect 22876 29260 22932 29262
rect 24444 30828 24500 30884
rect 25228 31724 25284 31780
rect 24668 30156 24724 30212
rect 24332 29986 24388 29988
rect 24332 29934 24334 29986
rect 24334 29934 24386 29986
rect 24386 29934 24388 29986
rect 24332 29932 24388 29934
rect 25788 31500 25844 31556
rect 25788 31218 25844 31220
rect 25788 31166 25790 31218
rect 25790 31166 25842 31218
rect 25842 31166 25844 31218
rect 25788 31164 25844 31166
rect 29372 41970 29428 41972
rect 29372 41918 29374 41970
rect 29374 41918 29426 41970
rect 29426 41918 29428 41970
rect 29372 41916 29428 41918
rect 29148 40236 29204 40292
rect 29708 44322 29764 44324
rect 29708 44270 29710 44322
rect 29710 44270 29762 44322
rect 29762 44270 29764 44322
rect 29708 44268 29764 44270
rect 29820 44210 29876 44212
rect 29820 44158 29822 44210
rect 29822 44158 29874 44210
rect 29874 44158 29876 44210
rect 29820 44156 29876 44158
rect 29596 43538 29652 43540
rect 29596 43486 29598 43538
rect 29598 43486 29650 43538
rect 29650 43486 29652 43538
rect 29596 43484 29652 43486
rect 29932 43762 29988 43764
rect 29932 43710 29934 43762
rect 29934 43710 29986 43762
rect 29986 43710 29988 43762
rect 29932 43708 29988 43710
rect 30156 45164 30212 45220
rect 30156 43708 30212 43764
rect 30044 43596 30100 43652
rect 29708 43036 29764 43092
rect 29596 42978 29652 42980
rect 29596 42926 29598 42978
rect 29598 42926 29650 42978
rect 29650 42926 29652 42978
rect 29596 42924 29652 42926
rect 29820 41970 29876 41972
rect 29820 41918 29822 41970
rect 29822 41918 29874 41970
rect 29874 41918 29876 41970
rect 29820 41916 29876 41918
rect 29708 40626 29764 40628
rect 29708 40574 29710 40626
rect 29710 40574 29762 40626
rect 29762 40574 29764 40626
rect 29708 40572 29764 40574
rect 29596 40460 29652 40516
rect 29820 40236 29876 40292
rect 29148 39618 29204 39620
rect 29148 39566 29150 39618
rect 29150 39566 29202 39618
rect 29202 39566 29204 39618
rect 29148 39564 29204 39566
rect 29260 39340 29316 39396
rect 29484 38834 29540 38836
rect 29484 38782 29486 38834
rect 29486 38782 29538 38834
rect 29538 38782 29540 38834
rect 29484 38780 29540 38782
rect 29036 38444 29092 38500
rect 29260 38556 29316 38612
rect 28588 38050 28644 38052
rect 28588 37998 28590 38050
rect 28590 37998 28642 38050
rect 28642 37998 28644 38050
rect 28588 37996 28644 37998
rect 28924 37772 28980 37828
rect 28476 37436 28532 37492
rect 28588 37324 28644 37380
rect 28924 37266 28980 37268
rect 28924 37214 28926 37266
rect 28926 37214 28978 37266
rect 28978 37214 28980 37266
rect 28924 37212 28980 37214
rect 29260 38050 29316 38052
rect 29260 37998 29262 38050
rect 29262 37998 29314 38050
rect 29314 37998 29316 38050
rect 29260 37996 29316 37998
rect 29260 37324 29316 37380
rect 29484 37996 29540 38052
rect 28140 36370 28196 36372
rect 28140 36318 28142 36370
rect 28142 36318 28194 36370
rect 28194 36318 28196 36370
rect 28140 36316 28196 36318
rect 28252 35980 28308 36036
rect 28364 35922 28420 35924
rect 28364 35870 28366 35922
rect 28366 35870 28418 35922
rect 28418 35870 28420 35922
rect 28364 35868 28420 35870
rect 28140 33516 28196 33572
rect 27020 33234 27076 33236
rect 27020 33182 27022 33234
rect 27022 33182 27074 33234
rect 27074 33182 27076 33234
rect 27020 33180 27076 33182
rect 26908 32620 26964 32676
rect 26124 31724 26180 31780
rect 29260 36876 29316 36932
rect 29148 36764 29204 36820
rect 28812 35980 28868 36036
rect 29708 37938 29764 37940
rect 29708 37886 29710 37938
rect 29710 37886 29762 37938
rect 29762 37886 29764 37938
rect 29708 37884 29764 37886
rect 30156 42700 30212 42756
rect 30380 45724 30436 45780
rect 30492 45388 30548 45444
rect 30380 43538 30436 43540
rect 30380 43486 30382 43538
rect 30382 43486 30434 43538
rect 30434 43486 30436 43538
rect 30380 43484 30436 43486
rect 30380 42754 30436 42756
rect 30380 42702 30382 42754
rect 30382 42702 30434 42754
rect 30434 42702 30436 42754
rect 30380 42700 30436 42702
rect 30828 46284 30884 46340
rect 30604 44322 30660 44324
rect 30604 44270 30606 44322
rect 30606 44270 30658 44322
rect 30658 44270 30660 44322
rect 30604 44268 30660 44270
rect 31052 48300 31108 48356
rect 31164 49308 31220 49364
rect 31612 48802 31668 48804
rect 31612 48750 31614 48802
rect 31614 48750 31666 48802
rect 31666 48750 31668 48802
rect 31612 48748 31668 48750
rect 31948 48972 32004 49028
rect 31052 48130 31108 48132
rect 31052 48078 31054 48130
rect 31054 48078 31106 48130
rect 31106 48078 31108 48130
rect 31052 48076 31108 48078
rect 31164 47628 31220 47684
rect 31388 47570 31444 47572
rect 31388 47518 31390 47570
rect 31390 47518 31442 47570
rect 31442 47518 31444 47570
rect 31388 47516 31444 47518
rect 31388 46620 31444 46676
rect 31500 45890 31556 45892
rect 31500 45838 31502 45890
rect 31502 45838 31554 45890
rect 31554 45838 31556 45890
rect 31500 45836 31556 45838
rect 31164 45106 31220 45108
rect 31164 45054 31166 45106
rect 31166 45054 31218 45106
rect 31218 45054 31220 45106
rect 31164 45052 31220 45054
rect 31388 44492 31444 44548
rect 31164 44380 31220 44436
rect 30940 44268 30996 44324
rect 30604 43596 30660 43652
rect 30716 43484 30772 43540
rect 30828 42924 30884 42980
rect 30604 42364 30660 42420
rect 30044 41356 30100 41412
rect 30604 41916 30660 41972
rect 30828 41916 30884 41972
rect 30828 40626 30884 40628
rect 30828 40574 30830 40626
rect 30830 40574 30882 40626
rect 30882 40574 30884 40626
rect 30828 40572 30884 40574
rect 30156 40236 30212 40292
rect 29932 39564 29988 39620
rect 30156 38162 30212 38164
rect 30156 38110 30158 38162
rect 30158 38110 30210 38162
rect 30210 38110 30212 38162
rect 30156 38108 30212 38110
rect 30156 37660 30212 37716
rect 29484 35980 29540 36036
rect 29596 37212 29652 37268
rect 29372 35868 29428 35924
rect 30716 37436 30772 37492
rect 29932 36258 29988 36260
rect 29932 36206 29934 36258
rect 29934 36206 29986 36258
rect 29986 36206 29988 36258
rect 29932 36204 29988 36206
rect 31052 43708 31108 43764
rect 31388 43708 31444 43764
rect 31276 42588 31332 42644
rect 31724 47682 31780 47684
rect 31724 47630 31726 47682
rect 31726 47630 31778 47682
rect 31778 47630 31780 47682
rect 31724 47628 31780 47630
rect 31948 48300 32004 48356
rect 32060 48130 32116 48132
rect 32060 48078 32062 48130
rect 32062 48078 32114 48130
rect 32114 48078 32116 48130
rect 32060 48076 32116 48078
rect 31724 47292 31780 47348
rect 32060 47180 32116 47236
rect 31724 45500 31780 45556
rect 31836 44322 31892 44324
rect 31836 44270 31838 44322
rect 31838 44270 31890 44322
rect 31890 44270 31892 44322
rect 31836 44268 31892 44270
rect 31612 43932 31668 43988
rect 32732 50428 32788 50484
rect 32620 50370 32676 50372
rect 32620 50318 32622 50370
rect 32622 50318 32674 50370
rect 32674 50318 32676 50370
rect 32620 50316 32676 50318
rect 32844 50316 32900 50372
rect 32508 50092 32564 50148
rect 32396 49922 32452 49924
rect 32396 49870 32398 49922
rect 32398 49870 32450 49922
rect 32450 49870 32452 49922
rect 32396 49868 32452 49870
rect 32396 48802 32452 48804
rect 32396 48750 32398 48802
rect 32398 48750 32450 48802
rect 32450 48750 32452 48802
rect 32396 48748 32452 48750
rect 33628 54684 33684 54740
rect 33628 54124 33684 54180
rect 35308 55970 35364 55972
rect 35308 55918 35310 55970
rect 35310 55918 35362 55970
rect 35362 55918 35364 55970
rect 35308 55916 35364 55918
rect 36092 55970 36148 55972
rect 36092 55918 36094 55970
rect 36094 55918 36146 55970
rect 36146 55918 36148 55970
rect 36092 55916 36148 55918
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 34860 55186 34916 55188
rect 34860 55134 34862 55186
rect 34862 55134 34914 55186
rect 34914 55134 34916 55186
rect 34860 55132 34916 55134
rect 34300 55020 34356 55076
rect 34748 54684 34804 54740
rect 33852 53452 33908 53508
rect 33628 53170 33684 53172
rect 33628 53118 33630 53170
rect 33630 53118 33682 53170
rect 33682 53118 33684 53170
rect 33628 53116 33684 53118
rect 33964 54348 34020 54404
rect 34076 53954 34132 53956
rect 34076 53902 34078 53954
rect 34078 53902 34130 53954
rect 34130 53902 34132 53954
rect 34076 53900 34132 53902
rect 34300 54124 34356 54180
rect 35980 55356 36036 55412
rect 34524 53564 34580 53620
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 35420 53900 35476 53956
rect 35196 53842 35252 53844
rect 35196 53790 35198 53842
rect 35198 53790 35250 53842
rect 35250 53790 35252 53842
rect 35196 53788 35252 53790
rect 34860 53116 34916 53172
rect 35420 53170 35476 53172
rect 35420 53118 35422 53170
rect 35422 53118 35474 53170
rect 35474 53118 35476 53170
rect 35420 53116 35476 53118
rect 34972 53058 35028 53060
rect 34972 53006 34974 53058
rect 34974 53006 35026 53058
rect 35026 53006 35028 53058
rect 34972 53004 35028 53006
rect 34524 52668 34580 52724
rect 33180 50988 33236 51044
rect 33292 51100 33348 51156
rect 33740 51548 33796 51604
rect 33516 50316 33572 50372
rect 33740 50594 33796 50596
rect 33740 50542 33742 50594
rect 33742 50542 33794 50594
rect 33794 50542 33796 50594
rect 33740 50540 33796 50542
rect 34188 50876 34244 50932
rect 34188 50540 34244 50596
rect 33404 49026 33460 49028
rect 33404 48974 33406 49026
rect 33406 48974 33458 49026
rect 33458 48974 33460 49026
rect 33404 48972 33460 48974
rect 32844 48076 32900 48132
rect 32956 48188 33012 48244
rect 32844 47740 32900 47796
rect 32172 46956 32228 47012
rect 32060 43148 32116 43204
rect 32396 47292 32452 47348
rect 32060 42924 32116 42980
rect 31836 42754 31892 42756
rect 31836 42702 31838 42754
rect 31838 42702 31890 42754
rect 31890 42702 31892 42754
rect 31836 42700 31892 42702
rect 31164 42530 31220 42532
rect 31164 42478 31166 42530
rect 31166 42478 31218 42530
rect 31218 42478 31220 42530
rect 31164 42476 31220 42478
rect 31164 42028 31220 42084
rect 31612 42530 31668 42532
rect 31612 42478 31614 42530
rect 31614 42478 31666 42530
rect 31666 42478 31668 42530
rect 31612 42476 31668 42478
rect 31500 41916 31556 41972
rect 31276 41356 31332 41412
rect 31388 41244 31444 41300
rect 31500 41186 31556 41188
rect 31500 41134 31502 41186
rect 31502 41134 31554 41186
rect 31554 41134 31556 41186
rect 31500 41132 31556 41134
rect 30940 38332 30996 38388
rect 31164 38050 31220 38052
rect 31164 37998 31166 38050
rect 31166 37998 31218 38050
rect 31218 37998 31220 38050
rect 31164 37996 31220 37998
rect 30156 36988 30212 37044
rect 30380 36652 30436 36708
rect 30716 36370 30772 36372
rect 30716 36318 30718 36370
rect 30718 36318 30770 36370
rect 30770 36318 30772 36370
rect 30716 36316 30772 36318
rect 29372 35698 29428 35700
rect 29372 35646 29374 35698
rect 29374 35646 29426 35698
rect 29426 35646 29428 35698
rect 29372 35644 29428 35646
rect 28700 34860 28756 34916
rect 29148 35084 29204 35140
rect 29484 35196 29540 35252
rect 29708 35644 29764 35700
rect 29484 34636 29540 34692
rect 30044 35196 30100 35252
rect 30268 35196 30324 35252
rect 30156 34524 30212 34580
rect 30380 34300 30436 34356
rect 30604 34636 30660 34692
rect 30492 34188 30548 34244
rect 32284 46060 32340 46116
rect 32956 46844 33012 46900
rect 32844 46114 32900 46116
rect 32844 46062 32846 46114
rect 32846 46062 32898 46114
rect 32898 46062 32900 46114
rect 32844 46060 32900 46062
rect 33516 47740 33572 47796
rect 33180 46898 33236 46900
rect 33180 46846 33182 46898
rect 33182 46846 33234 46898
rect 33234 46846 33236 46898
rect 33180 46844 33236 46846
rect 32508 45388 32564 45444
rect 32620 45612 32676 45668
rect 32508 45106 32564 45108
rect 32508 45054 32510 45106
rect 32510 45054 32562 45106
rect 32562 45054 32564 45106
rect 32508 45052 32564 45054
rect 32284 44492 32340 44548
rect 32732 44380 32788 44436
rect 32284 43820 32340 43876
rect 33068 44380 33124 44436
rect 33068 44210 33124 44212
rect 33068 44158 33070 44210
rect 33070 44158 33122 44210
rect 33122 44158 33124 44210
rect 33068 44156 33124 44158
rect 32844 43708 32900 43764
rect 33180 42924 33236 42980
rect 32396 42754 32452 42756
rect 32396 42702 32398 42754
rect 32398 42702 32450 42754
rect 32450 42702 32452 42754
rect 32396 42700 32452 42702
rect 32508 42642 32564 42644
rect 32508 42590 32510 42642
rect 32510 42590 32562 42642
rect 32562 42590 32564 42642
rect 32508 42588 32564 42590
rect 32732 42642 32788 42644
rect 32732 42590 32734 42642
rect 32734 42590 32786 42642
rect 32786 42590 32788 42642
rect 32732 42588 32788 42590
rect 32172 40796 32228 40852
rect 31500 40402 31556 40404
rect 31500 40350 31502 40402
rect 31502 40350 31554 40402
rect 31554 40350 31556 40402
rect 31500 40348 31556 40350
rect 31948 40348 32004 40404
rect 31724 40124 31780 40180
rect 32060 40124 32116 40180
rect 31948 39564 32004 39620
rect 31724 39228 31780 39284
rect 32060 39116 32116 39172
rect 32060 38668 32116 38724
rect 32284 39676 32340 39732
rect 32508 38722 32564 38724
rect 32508 38670 32510 38722
rect 32510 38670 32562 38722
rect 32562 38670 32564 38722
rect 32508 38668 32564 38670
rect 31276 37100 31332 37156
rect 31948 37212 32004 37268
rect 32172 37378 32228 37380
rect 32172 37326 32174 37378
rect 32174 37326 32226 37378
rect 32226 37326 32228 37378
rect 32172 37324 32228 37326
rect 32284 37212 32340 37268
rect 32844 38444 32900 38500
rect 32620 37660 32676 37716
rect 32060 36876 32116 36932
rect 31500 36540 31556 36596
rect 30940 36370 30996 36372
rect 30940 36318 30942 36370
rect 30942 36318 30994 36370
rect 30994 36318 30996 36370
rect 30940 36316 30996 36318
rect 31052 35196 31108 35252
rect 30940 34860 30996 34916
rect 32060 36316 32116 36372
rect 32172 37100 32228 37156
rect 32060 34972 32116 35028
rect 32396 36988 32452 37044
rect 33740 47516 33796 47572
rect 33628 47458 33684 47460
rect 33628 47406 33630 47458
rect 33630 47406 33682 47458
rect 33682 47406 33684 47458
rect 33628 47404 33684 47406
rect 33628 46956 33684 47012
rect 33404 45218 33460 45220
rect 33404 45166 33406 45218
rect 33406 45166 33458 45218
rect 33458 45166 33460 45218
rect 33404 45164 33460 45166
rect 33404 44716 33460 44772
rect 33404 44044 33460 44100
rect 33404 43596 33460 43652
rect 33852 46508 33908 46564
rect 33628 44044 33684 44100
rect 33404 43148 33460 43204
rect 33740 43372 33796 43428
rect 33852 45052 33908 45108
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 34860 52108 34916 52164
rect 35420 52162 35476 52164
rect 35420 52110 35422 52162
rect 35422 52110 35474 52162
rect 35474 52110 35476 52162
rect 35420 52108 35476 52110
rect 35196 51548 35252 51604
rect 34860 51490 34916 51492
rect 34860 51438 34862 51490
rect 34862 51438 34914 51490
rect 34914 51438 34916 51490
rect 34860 51436 34916 51438
rect 36204 53788 36260 53844
rect 36092 53564 36148 53620
rect 35980 53506 36036 53508
rect 35980 53454 35982 53506
rect 35982 53454 36034 53506
rect 36034 53454 36036 53506
rect 35980 53452 36036 53454
rect 35644 52332 35700 52388
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 35196 50652 35252 50708
rect 38556 57484 38612 57540
rect 37100 56700 37156 56756
rect 36988 56082 37044 56084
rect 36988 56030 36990 56082
rect 36990 56030 37042 56082
rect 37042 56030 37044 56082
rect 36988 56028 37044 56030
rect 36540 55468 36596 55524
rect 36428 55186 36484 55188
rect 36428 55134 36430 55186
rect 36430 55134 36482 55186
rect 36482 55134 36484 55186
rect 36428 55132 36484 55134
rect 36652 55020 36708 55076
rect 36988 54796 37044 54852
rect 36764 53788 36820 53844
rect 36428 52892 36484 52948
rect 36316 50428 36372 50484
rect 35420 49810 35476 49812
rect 35420 49758 35422 49810
rect 35422 49758 35474 49810
rect 35474 49758 35476 49810
rect 35420 49756 35476 49758
rect 34972 49698 35028 49700
rect 34972 49646 34974 49698
rect 34974 49646 35026 49698
rect 35026 49646 35028 49698
rect 34972 49644 35028 49646
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 34188 47346 34244 47348
rect 34188 47294 34190 47346
rect 34190 47294 34242 47346
rect 34242 47294 34244 47346
rect 34188 47292 34244 47294
rect 34076 46172 34132 46228
rect 34412 48972 34468 49028
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 35308 47516 35364 47572
rect 34300 45836 34356 45892
rect 34076 45218 34132 45220
rect 34076 45166 34078 45218
rect 34078 45166 34130 45218
rect 34130 45166 34132 45218
rect 34076 45164 34132 45166
rect 34300 44716 34356 44772
rect 33740 42194 33796 42196
rect 33740 42142 33742 42194
rect 33742 42142 33794 42194
rect 33794 42142 33796 42194
rect 33740 42140 33796 42142
rect 33628 41356 33684 41412
rect 33964 43708 34020 43764
rect 34188 43932 34244 43988
rect 34524 44940 34580 44996
rect 36316 49756 36372 49812
rect 35756 47682 35812 47684
rect 35756 47630 35758 47682
rect 35758 47630 35810 47682
rect 35810 47630 35812 47682
rect 35756 47628 35812 47630
rect 35532 46956 35588 47012
rect 35868 47292 35924 47348
rect 35980 47628 36036 47684
rect 36204 46620 36260 46676
rect 36876 53564 36932 53620
rect 36988 53116 37044 53172
rect 36988 52780 37044 52836
rect 36428 49138 36484 49140
rect 36428 49086 36430 49138
rect 36430 49086 36482 49138
rect 36482 49086 36484 49138
rect 36428 49084 36484 49086
rect 34748 44828 34804 44884
rect 34748 44380 34804 44436
rect 34524 43820 34580 43876
rect 34300 42924 34356 42980
rect 34188 41970 34244 41972
rect 34188 41918 34190 41970
rect 34190 41918 34242 41970
rect 34242 41918 34244 41970
rect 34188 41916 34244 41918
rect 34412 41468 34468 41524
rect 33852 40012 33908 40068
rect 34076 41020 34132 41076
rect 33516 39730 33572 39732
rect 33516 39678 33518 39730
rect 33518 39678 33570 39730
rect 33570 39678 33572 39730
rect 33516 39676 33572 39678
rect 33516 39116 33572 39172
rect 33404 39058 33460 39060
rect 33404 39006 33406 39058
rect 33406 39006 33458 39058
rect 33458 39006 33460 39058
rect 33404 39004 33460 39006
rect 33068 38050 33124 38052
rect 33068 37998 33070 38050
rect 33070 37998 33122 38050
rect 33122 37998 33124 38050
rect 33068 37996 33124 37998
rect 33292 38274 33348 38276
rect 33292 38222 33294 38274
rect 33294 38222 33346 38274
rect 33346 38222 33348 38274
rect 33292 38220 33348 38222
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 35308 45106 35364 45108
rect 35308 45054 35310 45106
rect 35310 45054 35362 45106
rect 35362 45054 35364 45106
rect 35308 45052 35364 45054
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 35084 44268 35140 44324
rect 35868 44268 35924 44324
rect 34860 43820 34916 43876
rect 34636 43650 34692 43652
rect 34636 43598 34638 43650
rect 34638 43598 34690 43650
rect 34690 43598 34692 43650
rect 34636 43596 34692 43598
rect 34860 43372 34916 43428
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 35532 42642 35588 42644
rect 35532 42590 35534 42642
rect 35534 42590 35586 42642
rect 35586 42590 35588 42642
rect 35532 42588 35588 42590
rect 35756 44098 35812 44100
rect 35756 44046 35758 44098
rect 35758 44046 35810 44098
rect 35810 44046 35812 44098
rect 35756 44044 35812 44046
rect 35644 42252 35700 42308
rect 34972 42140 35028 42196
rect 34860 42082 34916 42084
rect 34860 42030 34862 42082
rect 34862 42030 34914 42082
rect 34914 42030 34916 42082
rect 34860 42028 34916 42030
rect 35196 41970 35252 41972
rect 35196 41918 35198 41970
rect 35198 41918 35250 41970
rect 35250 41918 35252 41970
rect 35196 41916 35252 41918
rect 34972 41858 35028 41860
rect 34972 41806 34974 41858
rect 34974 41806 35026 41858
rect 35026 41806 35028 41858
rect 34972 41804 35028 41806
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 36428 44882 36484 44884
rect 36428 44830 36430 44882
rect 36430 44830 36482 44882
rect 36482 44830 36484 44882
rect 36428 44828 36484 44830
rect 36316 44098 36372 44100
rect 36316 44046 36318 44098
rect 36318 44046 36370 44098
rect 36370 44046 36372 44098
rect 36316 44044 36372 44046
rect 36652 49810 36708 49812
rect 36652 49758 36654 49810
rect 36654 49758 36706 49810
rect 36706 49758 36708 49810
rect 36652 49756 36708 49758
rect 37436 56194 37492 56196
rect 37436 56142 37438 56194
rect 37438 56142 37490 56194
rect 37490 56142 37492 56194
rect 37436 56140 37492 56142
rect 37884 55410 37940 55412
rect 37884 55358 37886 55410
rect 37886 55358 37938 55410
rect 37938 55358 37940 55410
rect 37884 55356 37940 55358
rect 37324 55074 37380 55076
rect 37324 55022 37326 55074
rect 37326 55022 37378 55074
rect 37378 55022 37380 55074
rect 37324 55020 37380 55022
rect 38220 55244 38276 55300
rect 37996 55074 38052 55076
rect 37996 55022 37998 55074
rect 37998 55022 38050 55074
rect 38050 55022 38052 55074
rect 37996 55020 38052 55022
rect 37212 53900 37268 53956
rect 38220 54684 38276 54740
rect 37660 54626 37716 54628
rect 37660 54574 37662 54626
rect 37662 54574 37714 54626
rect 37714 54574 37716 54626
rect 37660 54572 37716 54574
rect 38220 54514 38276 54516
rect 38220 54462 38222 54514
rect 38222 54462 38274 54514
rect 38274 54462 38276 54514
rect 38220 54460 38276 54462
rect 37324 51436 37380 51492
rect 37100 50988 37156 51044
rect 36988 50876 37044 50932
rect 37548 51884 37604 51940
rect 37436 50652 37492 50708
rect 40572 57372 40628 57428
rect 40460 57148 40516 57204
rect 40348 55298 40404 55300
rect 40348 55246 40350 55298
rect 40350 55246 40402 55298
rect 40402 55246 40404 55298
rect 40348 55244 40404 55246
rect 38780 55074 38836 55076
rect 38780 55022 38782 55074
rect 38782 55022 38834 55074
rect 38834 55022 38836 55074
rect 38780 55020 38836 55022
rect 38892 54402 38948 54404
rect 38892 54350 38894 54402
rect 38894 54350 38946 54402
rect 38946 54350 38948 54402
rect 38892 54348 38948 54350
rect 39004 53676 39060 53732
rect 37996 53170 38052 53172
rect 37996 53118 37998 53170
rect 37998 53118 38050 53170
rect 38050 53118 38052 53170
rect 37996 53116 38052 53118
rect 38444 53116 38500 53172
rect 39004 53506 39060 53508
rect 39004 53454 39006 53506
rect 39006 53454 39058 53506
rect 39058 53454 39060 53506
rect 39004 53452 39060 53454
rect 37996 52332 38052 52388
rect 36876 49532 36932 49588
rect 37772 50988 37828 51044
rect 36764 46956 36820 47012
rect 37324 49138 37380 49140
rect 37324 49086 37326 49138
rect 37326 49086 37378 49138
rect 37378 49086 37380 49138
rect 37324 49084 37380 49086
rect 38892 53004 38948 53060
rect 39788 54514 39844 54516
rect 39788 54462 39790 54514
rect 39790 54462 39842 54514
rect 39842 54462 39844 54514
rect 39788 54460 39844 54462
rect 39564 54402 39620 54404
rect 39564 54350 39566 54402
rect 39566 54350 39618 54402
rect 39618 54350 39620 54402
rect 39564 54348 39620 54350
rect 39788 53900 39844 53956
rect 39676 53452 39732 53508
rect 39004 52892 39060 52948
rect 39228 53004 39284 53060
rect 38444 51938 38500 51940
rect 38444 51886 38446 51938
rect 38446 51886 38498 51938
rect 38498 51886 38500 51938
rect 38444 51884 38500 51886
rect 38108 51436 38164 51492
rect 38108 50818 38164 50820
rect 38108 50766 38110 50818
rect 38110 50766 38162 50818
rect 38162 50766 38164 50818
rect 38108 50764 38164 50766
rect 38332 50652 38388 50708
rect 37996 50594 38052 50596
rect 37996 50542 37998 50594
rect 37998 50542 38050 50594
rect 38050 50542 38052 50594
rect 37996 50540 38052 50542
rect 38780 50428 38836 50484
rect 39564 53170 39620 53172
rect 39564 53118 39566 53170
rect 39566 53118 39618 53170
rect 39618 53118 39620 53170
rect 39564 53116 39620 53118
rect 40012 53842 40068 53844
rect 40012 53790 40014 53842
rect 40014 53790 40066 53842
rect 40066 53790 40068 53842
rect 40012 53788 40068 53790
rect 40348 53618 40404 53620
rect 40348 53566 40350 53618
rect 40350 53566 40402 53618
rect 40402 53566 40404 53618
rect 40348 53564 40404 53566
rect 40124 53170 40180 53172
rect 40124 53118 40126 53170
rect 40126 53118 40178 53170
rect 40178 53118 40180 53170
rect 40124 53116 40180 53118
rect 39452 53058 39508 53060
rect 39452 53006 39454 53058
rect 39454 53006 39506 53058
rect 39506 53006 39508 53058
rect 39452 53004 39508 53006
rect 40012 53004 40068 53060
rect 39452 52220 39508 52276
rect 39676 51938 39732 51940
rect 39676 51886 39678 51938
rect 39678 51886 39730 51938
rect 39730 51886 39732 51938
rect 39676 51884 39732 51886
rect 40236 52108 40292 52164
rect 39564 50652 39620 50708
rect 38444 49980 38500 50036
rect 37996 49084 38052 49140
rect 37100 48076 37156 48132
rect 37212 47458 37268 47460
rect 37212 47406 37214 47458
rect 37214 47406 37266 47458
rect 37266 47406 37268 47458
rect 37212 47404 37268 47406
rect 36988 46508 37044 46564
rect 36652 45724 36708 45780
rect 36876 45500 36932 45556
rect 36764 44156 36820 44212
rect 36428 43538 36484 43540
rect 36428 43486 36430 43538
rect 36430 43486 36482 43538
rect 36482 43486 36484 43538
rect 36428 43484 36484 43486
rect 36316 42978 36372 42980
rect 36316 42926 36318 42978
rect 36318 42926 36370 42978
rect 36370 42926 36372 42978
rect 36316 42924 36372 42926
rect 34748 41020 34804 41076
rect 35084 40402 35140 40404
rect 35084 40350 35086 40402
rect 35086 40350 35138 40402
rect 35138 40350 35140 40402
rect 35084 40348 35140 40350
rect 34300 39340 34356 39396
rect 34412 39564 34468 39620
rect 34188 38780 34244 38836
rect 34412 38668 34468 38724
rect 34188 38162 34244 38164
rect 34188 38110 34190 38162
rect 34190 38110 34242 38162
rect 34242 38110 34244 38162
rect 34188 38108 34244 38110
rect 33516 37548 33572 37604
rect 33180 37212 33236 37268
rect 33068 36876 33124 36932
rect 32956 36652 33012 36708
rect 34300 37826 34356 37828
rect 34300 37774 34302 37826
rect 34302 37774 34354 37826
rect 34354 37774 34356 37826
rect 34300 37772 34356 37774
rect 33964 36482 34020 36484
rect 33964 36430 33966 36482
rect 33966 36430 34018 36482
rect 34018 36430 34020 36482
rect 33964 36428 34020 36430
rect 34076 36370 34132 36372
rect 34076 36318 34078 36370
rect 34078 36318 34130 36370
rect 34130 36318 34132 36370
rect 34076 36316 34132 36318
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 36652 42588 36708 42644
rect 36652 42252 36708 42308
rect 36540 40962 36596 40964
rect 36540 40910 36542 40962
rect 36542 40910 36594 40962
rect 36594 40910 36596 40962
rect 36540 40908 36596 40910
rect 36092 39676 36148 39732
rect 34860 39618 34916 39620
rect 34860 39566 34862 39618
rect 34862 39566 34914 39618
rect 34914 39566 34916 39618
rect 34860 39564 34916 39566
rect 35756 39506 35812 39508
rect 35756 39454 35758 39506
rect 35758 39454 35810 39506
rect 35810 39454 35812 39506
rect 35756 39452 35812 39454
rect 35980 39394 36036 39396
rect 35980 39342 35982 39394
rect 35982 39342 36034 39394
rect 36034 39342 36036 39394
rect 35980 39340 36036 39342
rect 36316 39004 36372 39060
rect 34860 38946 34916 38948
rect 34860 38894 34862 38946
rect 34862 38894 34914 38946
rect 34914 38894 34916 38946
rect 34860 38892 34916 38894
rect 35756 38946 35812 38948
rect 35756 38894 35758 38946
rect 35758 38894 35810 38946
rect 35810 38894 35812 38946
rect 35756 38892 35812 38894
rect 34860 37324 34916 37380
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 32508 35420 32564 35476
rect 33852 36092 33908 36148
rect 33180 35420 33236 35476
rect 32060 34300 32116 34356
rect 28588 32732 28644 32788
rect 29484 32732 29540 32788
rect 29820 32786 29876 32788
rect 29820 32734 29822 32786
rect 29822 32734 29874 32786
rect 29874 32734 29876 32786
rect 29820 32732 29876 32734
rect 30156 32562 30212 32564
rect 30156 32510 30158 32562
rect 30158 32510 30210 32562
rect 30210 32510 30212 32562
rect 30156 32508 30212 32510
rect 29260 32396 29316 32452
rect 28476 31724 28532 31780
rect 25564 30828 25620 30884
rect 28140 31276 28196 31332
rect 26908 30994 26964 30996
rect 26908 30942 26910 30994
rect 26910 30942 26962 30994
rect 26962 30942 26964 30994
rect 26908 30940 26964 30942
rect 25900 30828 25956 30884
rect 26236 30882 26292 30884
rect 26236 30830 26238 30882
rect 26238 30830 26290 30882
rect 26290 30830 26292 30882
rect 26236 30828 26292 30830
rect 27804 30268 27860 30324
rect 25116 29596 25172 29652
rect 24668 29484 24724 29540
rect 25676 29932 25732 29988
rect 25452 29484 25508 29540
rect 26236 29538 26292 29540
rect 26236 29486 26238 29538
rect 26238 29486 26290 29538
rect 26290 29486 26292 29538
rect 26236 29484 26292 29486
rect 22540 27804 22596 27860
rect 22764 28642 22820 28644
rect 22764 28590 22766 28642
rect 22766 28590 22818 28642
rect 22818 28590 22820 28642
rect 22764 28588 22820 28590
rect 21532 25394 21588 25396
rect 21532 25342 21534 25394
rect 21534 25342 21586 25394
rect 21586 25342 21588 25394
rect 21532 25340 21588 25342
rect 21756 26236 21812 26292
rect 22204 25900 22260 25956
rect 20748 24050 20804 24052
rect 20748 23998 20750 24050
rect 20750 23998 20802 24050
rect 20802 23998 20804 24050
rect 20748 23996 20804 23998
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 20300 23100 20356 23156
rect 20188 22764 20244 22820
rect 19740 22370 19796 22372
rect 19740 22318 19742 22370
rect 19742 22318 19794 22370
rect 19794 22318 19796 22370
rect 19740 22316 19796 22318
rect 20188 22370 20244 22372
rect 20188 22318 20190 22370
rect 20190 22318 20242 22370
rect 20242 22318 20244 22370
rect 20188 22316 20244 22318
rect 20412 22316 20468 22372
rect 19292 21420 19348 21476
rect 19404 20802 19460 20804
rect 19404 20750 19406 20802
rect 19406 20750 19458 20802
rect 19458 20750 19460 20802
rect 19404 20748 19460 20750
rect 19068 19180 19124 19236
rect 19180 20188 19236 20244
rect 19404 20412 19460 20468
rect 19292 19740 19348 19796
rect 19292 19180 19348 19236
rect 19180 18956 19236 19012
rect 19068 18060 19124 18116
rect 19404 18674 19460 18676
rect 19404 18622 19406 18674
rect 19406 18622 19458 18674
rect 19458 18622 19460 18674
rect 19404 18620 19460 18622
rect 19292 17724 19348 17780
rect 18844 16268 18900 16324
rect 18732 15314 18788 15316
rect 18732 15262 18734 15314
rect 18734 15262 18786 15314
rect 18786 15262 18788 15314
rect 18732 15260 18788 15262
rect 18396 13634 18452 13636
rect 18396 13582 18398 13634
rect 18398 13582 18450 13634
rect 18450 13582 18452 13634
rect 18396 13580 18452 13582
rect 17500 12348 17556 12404
rect 17612 12796 17668 12852
rect 17500 11788 17556 11844
rect 17388 11394 17444 11396
rect 17388 11342 17390 11394
rect 17390 11342 17442 11394
rect 17442 11342 17444 11394
rect 17388 11340 17444 11342
rect 17276 9548 17332 9604
rect 16828 8988 16884 9044
rect 17164 8652 17220 8708
rect 16716 8316 16772 8372
rect 16828 8258 16884 8260
rect 16828 8206 16830 8258
rect 16830 8206 16882 8258
rect 16882 8206 16884 8258
rect 16828 8204 16884 8206
rect 16044 6636 16100 6692
rect 16492 6524 16548 6580
rect 16268 5906 16324 5908
rect 16268 5854 16270 5906
rect 16270 5854 16322 5906
rect 16322 5854 16324 5906
rect 16268 5852 16324 5854
rect 15708 5516 15764 5572
rect 14924 4898 14980 4900
rect 14924 4846 14926 4898
rect 14926 4846 14978 4898
rect 14978 4846 14980 4898
rect 14924 4844 14980 4846
rect 15260 4620 15316 4676
rect 16604 5740 16660 5796
rect 15820 4844 15876 4900
rect 16380 4844 16436 4900
rect 16604 5404 16660 5460
rect 16940 6076 16996 6132
rect 16828 5404 16884 5460
rect 16604 5068 16660 5124
rect 15820 4172 15876 4228
rect 16492 3836 16548 3892
rect 15820 3666 15876 3668
rect 15820 3614 15822 3666
rect 15822 3614 15874 3666
rect 15874 3614 15876 3666
rect 15820 3612 15876 3614
rect 13244 2716 13300 2772
rect 16940 4844 16996 4900
rect 16940 3948 16996 4004
rect 17836 12348 17892 12404
rect 18172 11228 18228 11284
rect 18172 10780 18228 10836
rect 18060 10668 18116 10724
rect 18060 10332 18116 10388
rect 18060 9772 18116 9828
rect 18172 9548 18228 9604
rect 17276 5852 17332 5908
rect 17276 5628 17332 5684
rect 17388 8092 17444 8148
rect 17612 8652 17668 8708
rect 17388 5516 17444 5572
rect 17612 7586 17668 7588
rect 17612 7534 17614 7586
rect 17614 7534 17666 7586
rect 17666 7534 17668 7586
rect 17612 7532 17668 7534
rect 17948 7644 18004 7700
rect 17948 7420 18004 7476
rect 18172 8764 18228 8820
rect 18508 13468 18564 13524
rect 18396 11506 18452 11508
rect 18396 11454 18398 11506
rect 18398 11454 18450 11506
rect 18450 11454 18452 11506
rect 18396 11452 18452 11454
rect 18956 13692 19012 13748
rect 18956 13468 19012 13524
rect 18956 12124 19012 12180
rect 18956 11900 19012 11956
rect 18620 11452 18676 11508
rect 18508 10892 18564 10948
rect 18396 10444 18452 10500
rect 18396 9714 18452 9716
rect 18396 9662 18398 9714
rect 18398 9662 18450 9714
rect 18450 9662 18452 9714
rect 18396 9660 18452 9662
rect 18620 9772 18676 9828
rect 18396 9436 18452 9492
rect 18620 9548 18676 9604
rect 18396 8652 18452 8708
rect 18508 8540 18564 8596
rect 18172 8204 18228 8260
rect 18172 7868 18228 7924
rect 18396 8092 18452 8148
rect 18060 6748 18116 6804
rect 18284 6748 18340 6804
rect 17836 6076 17892 6132
rect 17276 4844 17332 4900
rect 17612 4562 17668 4564
rect 17612 4510 17614 4562
rect 17614 4510 17666 4562
rect 17666 4510 17668 4562
rect 17612 4508 17668 4510
rect 18060 5740 18116 5796
rect 17836 5122 17892 5124
rect 17836 5070 17838 5122
rect 17838 5070 17890 5122
rect 17890 5070 17892 5122
rect 17836 5068 17892 5070
rect 19180 16492 19236 16548
rect 20188 22092 20244 22148
rect 19628 21980 19684 22036
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19964 21756 20020 21812
rect 20300 21586 20356 21588
rect 20300 21534 20302 21586
rect 20302 21534 20354 21586
rect 20354 21534 20356 21586
rect 20300 21532 20356 21534
rect 19964 21196 20020 21252
rect 19852 20524 19908 20580
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 20076 19740 20132 19796
rect 20748 22482 20804 22484
rect 20748 22430 20750 22482
rect 20750 22430 20802 22482
rect 20802 22430 20804 22482
rect 20748 22428 20804 22430
rect 22316 25506 22372 25508
rect 22316 25454 22318 25506
rect 22318 25454 22370 25506
rect 22370 25454 22372 25506
rect 22316 25452 22372 25454
rect 21756 25228 21812 25284
rect 22316 24892 22372 24948
rect 20972 24834 21028 24836
rect 20972 24782 20974 24834
rect 20974 24782 21026 24834
rect 21026 24782 21028 24834
rect 20972 24780 21028 24782
rect 21420 24780 21476 24836
rect 20636 20748 20692 20804
rect 20972 22540 21028 22596
rect 20412 20524 20468 20580
rect 20636 20578 20692 20580
rect 20636 20526 20638 20578
rect 20638 20526 20690 20578
rect 20690 20526 20692 20578
rect 20636 20524 20692 20526
rect 20412 20076 20468 20132
rect 20412 19180 20468 19236
rect 20412 19010 20468 19012
rect 20412 18958 20414 19010
rect 20414 18958 20466 19010
rect 20466 18958 20468 19010
rect 20412 18956 20468 18958
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19628 18396 19684 18452
rect 20188 18060 20244 18116
rect 19628 17724 19684 17780
rect 20412 17836 20468 17892
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19292 15372 19348 15428
rect 19404 16770 19460 16772
rect 19404 16718 19406 16770
rect 19406 16718 19458 16770
rect 19458 16718 19460 16770
rect 19404 16716 19460 16718
rect 19292 14252 19348 14308
rect 19180 13804 19236 13860
rect 19180 11788 19236 11844
rect 19068 10780 19124 10836
rect 18956 10610 19012 10612
rect 18956 10558 18958 10610
rect 18958 10558 19010 10610
rect 19010 10558 19012 10610
rect 18956 10556 19012 10558
rect 19852 16658 19908 16660
rect 19852 16606 19854 16658
rect 19854 16606 19906 16658
rect 19906 16606 19908 16658
rect 19852 16604 19908 16606
rect 19964 16268 20020 16324
rect 19740 16210 19796 16212
rect 19740 16158 19742 16210
rect 19742 16158 19794 16210
rect 19794 16158 19796 16210
rect 19740 16156 19796 16158
rect 20636 17276 20692 17332
rect 20524 16380 20580 16436
rect 20524 15820 20580 15876
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19516 14028 19572 14084
rect 19628 15484 19684 15540
rect 19740 15372 19796 15428
rect 20188 15036 20244 15092
rect 19740 14252 19796 14308
rect 20188 14812 20244 14868
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19740 13804 19796 13860
rect 20076 13522 20132 13524
rect 20076 13470 20078 13522
rect 20078 13470 20130 13522
rect 20130 13470 20132 13522
rect 20076 13468 20132 13470
rect 20188 13020 20244 13076
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19516 11228 19572 11284
rect 19404 10668 19460 10724
rect 19516 10610 19572 10612
rect 19516 10558 19518 10610
rect 19518 10558 19570 10610
rect 19570 10558 19572 10610
rect 19516 10556 19572 10558
rect 19292 10108 19348 10164
rect 21308 23714 21364 23716
rect 21308 23662 21310 23714
rect 21310 23662 21362 23714
rect 21362 23662 21364 23714
rect 21308 23660 21364 23662
rect 21196 22428 21252 22484
rect 21532 24556 21588 24612
rect 21868 24556 21924 24612
rect 21532 23996 21588 24052
rect 21084 21644 21140 21700
rect 21420 23154 21476 23156
rect 21420 23102 21422 23154
rect 21422 23102 21474 23154
rect 21474 23102 21476 23154
rect 21420 23100 21476 23102
rect 21420 22370 21476 22372
rect 21420 22318 21422 22370
rect 21422 22318 21474 22370
rect 21474 22318 21476 22370
rect 21420 22316 21476 22318
rect 21084 21084 21140 21140
rect 20860 19906 20916 19908
rect 20860 19854 20862 19906
rect 20862 19854 20914 19906
rect 20914 19854 20916 19906
rect 20860 19852 20916 19854
rect 20860 16882 20916 16884
rect 20860 16830 20862 16882
rect 20862 16830 20914 16882
rect 20914 16830 20916 16882
rect 20860 16828 20916 16830
rect 21756 24332 21812 24388
rect 21644 22092 21700 22148
rect 21532 21308 21588 21364
rect 21420 19740 21476 19796
rect 21308 18450 21364 18452
rect 21308 18398 21310 18450
rect 21310 18398 21362 18450
rect 21362 18398 21364 18450
rect 21308 18396 21364 18398
rect 21644 20412 21700 20468
rect 21420 17554 21476 17556
rect 21420 17502 21422 17554
rect 21422 17502 21474 17554
rect 21474 17502 21476 17554
rect 21420 17500 21476 17502
rect 21196 16940 21252 16996
rect 21420 15596 21476 15652
rect 21532 17276 21588 17332
rect 21308 15484 21364 15540
rect 21420 15426 21476 15428
rect 21420 15374 21422 15426
rect 21422 15374 21474 15426
rect 21474 15374 21476 15426
rect 21420 15372 21476 15374
rect 20748 15036 20804 15092
rect 21644 16268 21700 16324
rect 20748 14812 20804 14868
rect 20636 14642 20692 14644
rect 20636 14590 20638 14642
rect 20638 14590 20690 14642
rect 20690 14590 20692 14642
rect 20636 14588 20692 14590
rect 20636 13916 20692 13972
rect 20636 13692 20692 13748
rect 20188 11900 20244 11956
rect 20412 12236 20468 12292
rect 19852 11116 19908 11172
rect 20188 11170 20244 11172
rect 20188 11118 20190 11170
rect 20190 11118 20242 11170
rect 20242 11118 20244 11170
rect 20188 11116 20244 11118
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19740 10780 19796 10836
rect 18732 9324 18788 9380
rect 18844 9436 18900 9492
rect 18732 8428 18788 8484
rect 18956 9266 19012 9268
rect 18956 9214 18958 9266
rect 18958 9214 19010 9266
rect 19010 9214 19012 9266
rect 18956 9212 19012 9214
rect 19292 9772 19348 9828
rect 19628 9714 19684 9716
rect 19628 9662 19630 9714
rect 19630 9662 19682 9714
rect 19682 9662 19684 9714
rect 19628 9660 19684 9662
rect 19180 9548 19236 9604
rect 19404 9602 19460 9604
rect 19404 9550 19406 9602
rect 19406 9550 19458 9602
rect 19458 9550 19460 9602
rect 19404 9548 19460 9550
rect 19740 9548 19796 9604
rect 19964 9884 20020 9940
rect 20300 10108 20356 10164
rect 19964 9548 20020 9604
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19068 9042 19124 9044
rect 19068 8990 19070 9042
rect 19070 8990 19122 9042
rect 19122 8990 19124 9042
rect 19068 8988 19124 8990
rect 19404 8876 19460 8932
rect 19180 8428 19236 8484
rect 18620 7474 18676 7476
rect 18620 7422 18622 7474
rect 18622 7422 18674 7474
rect 18674 7422 18676 7474
rect 18620 7420 18676 7422
rect 18508 7362 18564 7364
rect 18508 7310 18510 7362
rect 18510 7310 18562 7362
rect 18562 7310 18564 7362
rect 18508 7308 18564 7310
rect 18396 6690 18452 6692
rect 18396 6638 18398 6690
rect 18398 6638 18450 6690
rect 18450 6638 18452 6690
rect 18396 6636 18452 6638
rect 18732 7196 18788 7252
rect 18732 6524 18788 6580
rect 19068 6524 19124 6580
rect 18508 6412 18564 6468
rect 18508 5906 18564 5908
rect 18508 5854 18510 5906
rect 18510 5854 18562 5906
rect 18562 5854 18564 5906
rect 18508 5852 18564 5854
rect 18284 5292 18340 5348
rect 18396 5180 18452 5236
rect 18620 5122 18676 5124
rect 18620 5070 18622 5122
rect 18622 5070 18674 5122
rect 18674 5070 18676 5122
rect 18620 5068 18676 5070
rect 18956 6130 19012 6132
rect 18956 6078 18958 6130
rect 18958 6078 19010 6130
rect 19010 6078 19012 6130
rect 18956 6076 19012 6078
rect 18732 4956 18788 5012
rect 19628 8428 19684 8484
rect 20188 8764 20244 8820
rect 20188 8428 20244 8484
rect 19964 8146 20020 8148
rect 19964 8094 19966 8146
rect 19966 8094 20018 8146
rect 20018 8094 20020 8146
rect 19964 8092 20020 8094
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 20076 7698 20132 7700
rect 20076 7646 20078 7698
rect 20078 7646 20130 7698
rect 20130 7646 20132 7698
rect 20076 7644 20132 7646
rect 19964 7532 20020 7588
rect 21084 15036 21140 15092
rect 21084 14364 21140 14420
rect 21196 14476 21252 14532
rect 20972 13746 21028 13748
rect 20972 13694 20974 13746
rect 20974 13694 21026 13746
rect 21026 13694 21028 13746
rect 20972 13692 21028 13694
rect 20748 12908 20804 12964
rect 20860 11788 20916 11844
rect 20748 11676 20804 11732
rect 20524 10556 20580 10612
rect 20748 9996 20804 10052
rect 20636 9826 20692 9828
rect 20636 9774 20638 9826
rect 20638 9774 20690 9826
rect 20690 9774 20692 9826
rect 20636 9772 20692 9774
rect 20412 7644 20468 7700
rect 20524 9660 20580 9716
rect 20748 9602 20804 9604
rect 20748 9550 20750 9602
rect 20750 9550 20802 9602
rect 20802 9550 20804 9602
rect 20748 9548 20804 9550
rect 20524 8876 20580 8932
rect 20300 7420 20356 7476
rect 19404 7362 19460 7364
rect 19404 7310 19406 7362
rect 19406 7310 19458 7362
rect 19458 7310 19460 7362
rect 19404 7308 19460 7310
rect 19292 7196 19348 7252
rect 19628 6972 19684 7028
rect 19516 5906 19572 5908
rect 19516 5854 19518 5906
rect 19518 5854 19570 5906
rect 19570 5854 19572 5906
rect 19516 5852 19572 5854
rect 19852 6578 19908 6580
rect 19852 6526 19854 6578
rect 19854 6526 19906 6578
rect 19906 6526 19908 6578
rect 19852 6524 19908 6526
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 20188 6130 20244 6132
rect 20188 6078 20190 6130
rect 20190 6078 20242 6130
rect 20242 6078 20244 6130
rect 20188 6076 20244 6078
rect 19852 6018 19908 6020
rect 19852 5966 19854 6018
rect 19854 5966 19906 6018
rect 19906 5966 19908 6018
rect 19852 5964 19908 5966
rect 21084 11116 21140 11172
rect 21084 10332 21140 10388
rect 21532 14530 21588 14532
rect 21532 14478 21534 14530
rect 21534 14478 21586 14530
rect 21586 14478 21588 14530
rect 21532 14476 21588 14478
rect 21308 14140 21364 14196
rect 21532 13916 21588 13972
rect 21308 12178 21364 12180
rect 21308 12126 21310 12178
rect 21310 12126 21362 12178
rect 21362 12126 21364 12178
rect 21308 12124 21364 12126
rect 22092 24108 22148 24164
rect 21868 23548 21924 23604
rect 22540 25228 22596 25284
rect 22428 23324 22484 23380
rect 23100 28364 23156 28420
rect 22764 28028 22820 28084
rect 22764 27186 22820 27188
rect 22764 27134 22766 27186
rect 22766 27134 22818 27186
rect 22818 27134 22820 27186
rect 22764 27132 22820 27134
rect 22988 26460 23044 26516
rect 22316 22316 22372 22372
rect 22428 21532 22484 21588
rect 21868 21420 21924 21476
rect 22428 20300 22484 20356
rect 22540 20524 22596 20580
rect 21868 18620 21924 18676
rect 22428 20130 22484 20132
rect 22428 20078 22430 20130
rect 22430 20078 22482 20130
rect 22482 20078 22484 20130
rect 22428 20076 22484 20078
rect 22316 19292 22372 19348
rect 22316 19122 22372 19124
rect 22316 19070 22318 19122
rect 22318 19070 22370 19122
rect 22370 19070 22372 19122
rect 22316 19068 22372 19070
rect 24668 28530 24724 28532
rect 24668 28478 24670 28530
rect 24670 28478 24722 28530
rect 24722 28478 24724 28530
rect 24668 28476 24724 28478
rect 24668 28082 24724 28084
rect 24668 28030 24670 28082
rect 24670 28030 24722 28082
rect 24722 28030 24724 28082
rect 24668 28028 24724 28030
rect 23548 27468 23604 27524
rect 23212 25506 23268 25508
rect 23212 25454 23214 25506
rect 23214 25454 23266 25506
rect 23266 25454 23268 25506
rect 23212 25452 23268 25454
rect 23324 26908 23380 26964
rect 23212 24892 23268 24948
rect 23436 25900 23492 25956
rect 23324 24610 23380 24612
rect 23324 24558 23326 24610
rect 23326 24558 23378 24610
rect 23378 24558 23380 24610
rect 23324 24556 23380 24558
rect 23212 24444 23268 24500
rect 22988 23436 23044 23492
rect 22764 23042 22820 23044
rect 22764 22990 22766 23042
rect 22766 22990 22818 23042
rect 22818 22990 22820 23042
rect 22764 22988 22820 22990
rect 22764 20412 22820 20468
rect 22988 22540 23044 22596
rect 22988 22204 23044 22260
rect 23100 21586 23156 21588
rect 23100 21534 23102 21586
rect 23102 21534 23154 21586
rect 23154 21534 23156 21586
rect 23100 21532 23156 21534
rect 22540 18844 22596 18900
rect 22988 19404 23044 19460
rect 22428 18450 22484 18452
rect 22428 18398 22430 18450
rect 22430 18398 22482 18450
rect 22482 18398 22484 18450
rect 22428 18396 22484 18398
rect 22540 18172 22596 18228
rect 21868 16492 21924 16548
rect 21980 17612 22036 17668
rect 21980 15932 22036 15988
rect 22092 15820 22148 15876
rect 21980 15708 22036 15764
rect 21756 14812 21812 14868
rect 22876 19180 22932 19236
rect 21868 13580 21924 13636
rect 21756 12124 21812 12180
rect 21980 12572 22036 12628
rect 22316 16156 22372 16212
rect 21980 11900 22036 11956
rect 21868 11788 21924 11844
rect 22428 16098 22484 16100
rect 22428 16046 22430 16098
rect 22430 16046 22482 16098
rect 22482 16046 22484 16098
rect 22428 16044 22484 16046
rect 22764 16044 22820 16100
rect 22316 14364 22372 14420
rect 22204 14028 22260 14084
rect 21756 11004 21812 11060
rect 21084 9660 21140 9716
rect 21084 8540 21140 8596
rect 20972 7756 21028 7812
rect 20636 7644 20692 7700
rect 20748 6748 20804 6804
rect 20860 6860 20916 6916
rect 20524 6636 20580 6692
rect 20636 6466 20692 6468
rect 20636 6414 20638 6466
rect 20638 6414 20690 6466
rect 20690 6414 20692 6466
rect 20636 6412 20692 6414
rect 20412 5852 20468 5908
rect 18396 4562 18452 4564
rect 18396 4510 18398 4562
rect 18398 4510 18450 4562
rect 18450 4510 18452 4562
rect 18396 4508 18452 4510
rect 18284 4396 18340 4452
rect 18844 4450 18900 4452
rect 18844 4398 18846 4450
rect 18846 4398 18898 4450
rect 18898 4398 18900 4450
rect 18844 4396 18900 4398
rect 19852 5628 19908 5684
rect 19740 5292 19796 5348
rect 19292 4844 19348 4900
rect 19516 5180 19572 5236
rect 19180 4620 19236 4676
rect 19292 4450 19348 4452
rect 19292 4398 19294 4450
rect 19294 4398 19346 4450
rect 19346 4398 19348 4450
rect 19292 4396 19348 4398
rect 18620 4284 18676 4340
rect 19516 4844 19572 4900
rect 20524 5740 20580 5796
rect 20076 5180 20132 5236
rect 20300 5516 20356 5572
rect 20188 4898 20244 4900
rect 20188 4846 20190 4898
rect 20190 4846 20242 4898
rect 20242 4846 20244 4898
rect 20188 4844 20244 4846
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 19964 4562 20020 4564
rect 19964 4510 19966 4562
rect 19966 4510 20018 4562
rect 20018 4510 20020 4562
rect 19964 4508 20020 4510
rect 19292 3836 19348 3892
rect 19180 3612 19236 3668
rect 20524 5404 20580 5460
rect 20860 5628 20916 5684
rect 21084 6300 21140 6356
rect 21084 5516 21140 5572
rect 21196 6748 21252 6804
rect 20748 5292 20804 5348
rect 20636 5180 20692 5236
rect 21420 8370 21476 8372
rect 21420 8318 21422 8370
rect 21422 8318 21474 8370
rect 21474 8318 21476 8370
rect 21420 8316 21476 8318
rect 21644 9996 21700 10052
rect 21756 9938 21812 9940
rect 21756 9886 21758 9938
rect 21758 9886 21810 9938
rect 21810 9886 21812 9938
rect 21756 9884 21812 9886
rect 21980 9548 22036 9604
rect 22092 10108 22148 10164
rect 21644 8876 21700 8932
rect 21980 8428 22036 8484
rect 21532 8092 21588 8148
rect 21868 7698 21924 7700
rect 21868 7646 21870 7698
rect 21870 7646 21922 7698
rect 21922 7646 21924 7698
rect 21868 7644 21924 7646
rect 21644 7474 21700 7476
rect 21644 7422 21646 7474
rect 21646 7422 21698 7474
rect 21698 7422 21700 7474
rect 21644 7420 21700 7422
rect 21980 7196 22036 7252
rect 21756 6972 21812 7028
rect 21420 6690 21476 6692
rect 21420 6638 21422 6690
rect 21422 6638 21474 6690
rect 21474 6638 21476 6690
rect 21420 6636 21476 6638
rect 21644 6524 21700 6580
rect 21644 5906 21700 5908
rect 21644 5854 21646 5906
rect 21646 5854 21698 5906
rect 21698 5854 21700 5906
rect 21644 5852 21700 5854
rect 21532 5740 21588 5796
rect 20524 4060 20580 4116
rect 21308 5628 21364 5684
rect 22540 15596 22596 15652
rect 22764 15426 22820 15428
rect 22764 15374 22766 15426
rect 22766 15374 22818 15426
rect 22818 15374 22820 15426
rect 22764 15372 22820 15374
rect 22764 15202 22820 15204
rect 22764 15150 22766 15202
rect 22766 15150 22818 15202
rect 22818 15150 22820 15202
rect 22764 15148 22820 15150
rect 22652 14924 22708 14980
rect 22428 13804 22484 13860
rect 22428 12962 22484 12964
rect 22428 12910 22430 12962
rect 22430 12910 22482 12962
rect 22482 12910 22484 12962
rect 22428 12908 22484 12910
rect 22764 14700 22820 14756
rect 22988 18396 23044 18452
rect 23996 26012 24052 26068
rect 23884 25506 23940 25508
rect 23884 25454 23886 25506
rect 23886 25454 23938 25506
rect 23938 25454 23940 25506
rect 23884 25452 23940 25454
rect 23772 24108 23828 24164
rect 23996 23884 24052 23940
rect 25676 28028 25732 28084
rect 24332 26796 24388 26852
rect 24780 26348 24836 26404
rect 24332 26124 24388 26180
rect 23436 23436 23492 23492
rect 23324 22652 23380 22708
rect 24444 23436 24500 23492
rect 23436 22316 23492 22372
rect 23548 21644 23604 21700
rect 23436 21586 23492 21588
rect 23436 21534 23438 21586
rect 23438 21534 23490 21586
rect 23490 21534 23492 21586
rect 23436 21532 23492 21534
rect 24332 21756 24388 21812
rect 23884 21474 23940 21476
rect 23884 21422 23886 21474
rect 23886 21422 23938 21474
rect 23938 21422 23940 21474
rect 23884 21420 23940 21422
rect 24220 21362 24276 21364
rect 24220 21310 24222 21362
rect 24222 21310 24274 21362
rect 24274 21310 24276 21362
rect 24220 21308 24276 21310
rect 23436 20018 23492 20020
rect 23436 19966 23438 20018
rect 23438 19966 23490 20018
rect 23490 19966 23492 20018
rect 23436 19964 23492 19966
rect 24220 20130 24276 20132
rect 24220 20078 24222 20130
rect 24222 20078 24274 20130
rect 24274 20078 24276 20130
rect 24220 20076 24276 20078
rect 23996 19516 24052 19572
rect 24220 19516 24276 19572
rect 23884 19068 23940 19124
rect 23324 18844 23380 18900
rect 23324 18338 23380 18340
rect 23324 18286 23326 18338
rect 23326 18286 23378 18338
rect 23378 18286 23380 18338
rect 23324 18284 23380 18286
rect 23324 17836 23380 17892
rect 23772 18508 23828 18564
rect 23772 18226 23828 18228
rect 23772 18174 23774 18226
rect 23774 18174 23826 18226
rect 23826 18174 23828 18226
rect 23772 18172 23828 18174
rect 23772 17948 23828 18004
rect 23772 17778 23828 17780
rect 23772 17726 23774 17778
rect 23774 17726 23826 17778
rect 23826 17726 23828 17778
rect 23772 17724 23828 17726
rect 23548 17612 23604 17668
rect 22988 17500 23044 17556
rect 23100 16828 23156 16884
rect 23772 16994 23828 16996
rect 23772 16942 23774 16994
rect 23774 16942 23826 16994
rect 23826 16942 23828 16994
rect 23772 16940 23828 16942
rect 23436 16210 23492 16212
rect 23436 16158 23438 16210
rect 23438 16158 23490 16210
rect 23490 16158 23492 16210
rect 23436 16156 23492 16158
rect 23324 16098 23380 16100
rect 23324 16046 23326 16098
rect 23326 16046 23378 16098
rect 23378 16046 23380 16098
rect 23324 16044 23380 16046
rect 24668 25228 24724 25284
rect 24668 23100 24724 23156
rect 24892 22146 24948 22148
rect 24892 22094 24894 22146
rect 24894 22094 24946 22146
rect 24946 22094 24948 22146
rect 24892 22092 24948 22094
rect 24556 20524 24612 20580
rect 24332 17666 24388 17668
rect 24332 17614 24334 17666
rect 24334 17614 24386 17666
rect 24386 17614 24388 17666
rect 24332 17612 24388 17614
rect 24220 17388 24276 17444
rect 24332 17052 24388 17108
rect 25228 25788 25284 25844
rect 25116 25506 25172 25508
rect 25116 25454 25118 25506
rect 25118 25454 25170 25506
rect 25170 25454 25172 25506
rect 25116 25452 25172 25454
rect 25340 25228 25396 25284
rect 25452 27468 25508 27524
rect 25228 24892 25284 24948
rect 25340 24668 25396 24724
rect 25788 26962 25844 26964
rect 25788 26910 25790 26962
rect 25790 26910 25842 26962
rect 25842 26910 25844 26962
rect 25788 26908 25844 26910
rect 25788 26012 25844 26068
rect 25564 24722 25620 24724
rect 25564 24670 25566 24722
rect 25566 24670 25618 24722
rect 25618 24670 25620 24722
rect 25564 24668 25620 24670
rect 26124 28642 26180 28644
rect 26124 28590 26126 28642
rect 26126 28590 26178 28642
rect 26178 28590 26180 28642
rect 26124 28588 26180 28590
rect 26124 28028 26180 28084
rect 26908 28082 26964 28084
rect 26908 28030 26910 28082
rect 26910 28030 26962 28082
rect 26962 28030 26964 28082
rect 26908 28028 26964 28030
rect 27692 28082 27748 28084
rect 27692 28030 27694 28082
rect 27694 28030 27746 28082
rect 27746 28030 27748 28082
rect 27692 28028 27748 28030
rect 27468 27804 27524 27860
rect 26236 27132 26292 27188
rect 26460 27020 26516 27076
rect 27132 27020 27188 27076
rect 27244 26796 27300 26852
rect 26012 25900 26068 25956
rect 27356 26012 27412 26068
rect 26124 25340 26180 25396
rect 26572 24556 26628 24612
rect 25452 23714 25508 23716
rect 25452 23662 25454 23714
rect 25454 23662 25506 23714
rect 25506 23662 25508 23714
rect 25452 23660 25508 23662
rect 25340 23042 25396 23044
rect 25340 22990 25342 23042
rect 25342 22990 25394 23042
rect 25394 22990 25396 23042
rect 25340 22988 25396 22990
rect 25564 23436 25620 23492
rect 25340 21586 25396 21588
rect 25340 21534 25342 21586
rect 25342 21534 25394 21586
rect 25394 21534 25396 21586
rect 25340 21532 25396 21534
rect 25228 20972 25284 21028
rect 25340 20802 25396 20804
rect 25340 20750 25342 20802
rect 25342 20750 25394 20802
rect 25394 20750 25396 20802
rect 25340 20748 25396 20750
rect 25228 19964 25284 20020
rect 25340 20188 25396 20244
rect 25676 23154 25732 23156
rect 25676 23102 25678 23154
rect 25678 23102 25730 23154
rect 25730 23102 25732 23154
rect 25676 23100 25732 23102
rect 26460 23324 26516 23380
rect 26908 24610 26964 24612
rect 26908 24558 26910 24610
rect 26910 24558 26962 24610
rect 26962 24558 26964 24610
rect 26908 24556 26964 24558
rect 26684 23212 26740 23268
rect 26572 22764 26628 22820
rect 26572 22594 26628 22596
rect 26572 22542 26574 22594
rect 26574 22542 26626 22594
rect 26626 22542 26628 22594
rect 26572 22540 26628 22542
rect 26460 22370 26516 22372
rect 26460 22318 26462 22370
rect 26462 22318 26514 22370
rect 26514 22318 26516 22370
rect 26460 22316 26516 22318
rect 26684 22370 26740 22372
rect 26684 22318 26686 22370
rect 26686 22318 26738 22370
rect 26738 22318 26740 22370
rect 26684 22316 26740 22318
rect 26908 22652 26964 22708
rect 27020 22370 27076 22372
rect 27020 22318 27022 22370
rect 27022 22318 27074 22370
rect 27074 22318 27076 22370
rect 27020 22316 27076 22318
rect 25900 21868 25956 21924
rect 26012 21810 26068 21812
rect 26012 21758 26014 21810
rect 26014 21758 26066 21810
rect 26066 21758 26068 21810
rect 26012 21756 26068 21758
rect 26236 21698 26292 21700
rect 26236 21646 26238 21698
rect 26238 21646 26290 21698
rect 26290 21646 26292 21698
rect 26236 21644 26292 21646
rect 25676 20860 25732 20916
rect 25452 19740 25508 19796
rect 25116 19346 25172 19348
rect 25116 19294 25118 19346
rect 25118 19294 25170 19346
rect 25170 19294 25172 19346
rect 25116 19292 25172 19294
rect 24556 18284 24612 18340
rect 24556 17052 24612 17108
rect 23884 16044 23940 16100
rect 23996 15820 24052 15876
rect 24444 15820 24500 15876
rect 24444 15484 24500 15540
rect 23548 15036 23604 15092
rect 24108 14700 24164 14756
rect 23100 14364 23156 14420
rect 23660 14364 23716 14420
rect 23324 13916 23380 13972
rect 22988 13746 23044 13748
rect 22988 13694 22990 13746
rect 22990 13694 23042 13746
rect 23042 13694 23044 13746
rect 22988 13692 23044 13694
rect 22764 13468 22820 13524
rect 22764 13244 22820 13300
rect 23100 13244 23156 13300
rect 22428 12124 22484 12180
rect 22652 12124 22708 12180
rect 22652 11900 22708 11956
rect 22876 11900 22932 11956
rect 22540 11564 22596 11620
rect 22988 11564 23044 11620
rect 23212 12124 23268 12180
rect 22540 10722 22596 10724
rect 22540 10670 22542 10722
rect 22542 10670 22594 10722
rect 22594 10670 22596 10722
rect 22540 10668 22596 10670
rect 22764 10332 22820 10388
rect 22540 9714 22596 9716
rect 22540 9662 22542 9714
rect 22542 9662 22594 9714
rect 22594 9662 22596 9714
rect 22540 9660 22596 9662
rect 22652 9602 22708 9604
rect 22652 9550 22654 9602
rect 22654 9550 22706 9602
rect 22706 9550 22708 9602
rect 22652 9548 22708 9550
rect 22428 9436 22484 9492
rect 22764 9436 22820 9492
rect 22316 8428 22372 8484
rect 22428 8540 22484 8596
rect 23100 11394 23156 11396
rect 23100 11342 23102 11394
rect 23102 11342 23154 11394
rect 23154 11342 23156 11394
rect 23100 11340 23156 11342
rect 22988 10834 23044 10836
rect 22988 10782 22990 10834
rect 22990 10782 23042 10834
rect 23042 10782 23044 10834
rect 22988 10780 23044 10782
rect 22876 7868 22932 7924
rect 23100 10332 23156 10388
rect 23548 13916 23604 13972
rect 23548 13468 23604 13524
rect 23436 11564 23492 11620
rect 23772 13804 23828 13860
rect 23884 13244 23940 13300
rect 23772 11788 23828 11844
rect 23772 11394 23828 11396
rect 23772 11342 23774 11394
rect 23774 11342 23826 11394
rect 23826 11342 23828 11394
rect 23772 11340 23828 11342
rect 23884 11116 23940 11172
rect 23436 10108 23492 10164
rect 23324 9996 23380 10052
rect 23772 10668 23828 10724
rect 23324 8876 23380 8932
rect 23100 8764 23156 8820
rect 22204 6972 22260 7028
rect 22092 6636 22148 6692
rect 22316 5852 22372 5908
rect 21420 4508 21476 4564
rect 22204 5122 22260 5124
rect 22204 5070 22206 5122
rect 22206 5070 22258 5122
rect 22258 5070 22260 5122
rect 22204 5068 22260 5070
rect 22428 6412 22484 6468
rect 21868 4562 21924 4564
rect 21868 4510 21870 4562
rect 21870 4510 21922 4562
rect 21922 4510 21924 4562
rect 21868 4508 21924 4510
rect 21532 4396 21588 4452
rect 22204 4450 22260 4452
rect 22204 4398 22206 4450
rect 22206 4398 22258 4450
rect 22258 4398 22260 4450
rect 22204 4396 22260 4398
rect 21532 3948 21588 4004
rect 22652 6018 22708 6020
rect 22652 5966 22654 6018
rect 22654 5966 22706 6018
rect 22706 5966 22708 6018
rect 22652 5964 22708 5966
rect 22988 5906 23044 5908
rect 22988 5854 22990 5906
rect 22990 5854 23042 5906
rect 23042 5854 23044 5906
rect 22988 5852 23044 5854
rect 23100 5628 23156 5684
rect 23324 8428 23380 8484
rect 23212 5068 23268 5124
rect 23772 9436 23828 9492
rect 23884 9100 23940 9156
rect 24220 13020 24276 13076
rect 24444 12460 24500 12516
rect 24108 11340 24164 11396
rect 24220 11900 24276 11956
rect 25004 18620 25060 18676
rect 25228 19010 25284 19012
rect 25228 18958 25230 19010
rect 25230 18958 25282 19010
rect 25282 18958 25284 19010
rect 25228 18956 25284 18958
rect 26236 21084 26292 21140
rect 26012 20690 26068 20692
rect 26012 20638 26014 20690
rect 26014 20638 26066 20690
rect 26066 20638 26068 20690
rect 26012 20636 26068 20638
rect 26012 19906 26068 19908
rect 26012 19854 26014 19906
rect 26014 19854 26066 19906
rect 26066 19854 26068 19906
rect 26012 19852 26068 19854
rect 25788 19740 25844 19796
rect 25676 19516 25732 19572
rect 25452 18956 25508 19012
rect 26012 19234 26068 19236
rect 26012 19182 26014 19234
rect 26014 19182 26066 19234
rect 26066 19182 26068 19234
rect 26012 19180 26068 19182
rect 25564 18172 25620 18228
rect 25004 18060 25060 18116
rect 24668 16940 24724 16996
rect 25452 17724 25508 17780
rect 25340 16268 25396 16324
rect 25004 16098 25060 16100
rect 25004 16046 25006 16098
rect 25006 16046 25058 16098
rect 25058 16046 25060 16098
rect 25004 16044 25060 16046
rect 25116 15820 25172 15876
rect 24668 15426 24724 15428
rect 24668 15374 24670 15426
rect 24670 15374 24722 15426
rect 24722 15374 24724 15426
rect 24668 15372 24724 15374
rect 24892 15148 24948 15204
rect 24780 13804 24836 13860
rect 25116 14812 25172 14868
rect 25004 14252 25060 14308
rect 25564 16156 25620 16212
rect 25900 18284 25956 18340
rect 25900 17724 25956 17780
rect 26012 17612 26068 17668
rect 25788 16940 25844 16996
rect 25788 15596 25844 15652
rect 25676 15202 25732 15204
rect 25676 15150 25678 15202
rect 25678 15150 25730 15202
rect 25730 15150 25732 15202
rect 25676 15148 25732 15150
rect 25676 14700 25732 14756
rect 24332 11676 24388 11732
rect 24556 11900 24612 11956
rect 24892 11676 24948 11732
rect 25116 13186 25172 13188
rect 25116 13134 25118 13186
rect 25118 13134 25170 13186
rect 25170 13134 25172 13186
rect 25116 13132 25172 13134
rect 25004 11564 25060 11620
rect 25116 11788 25172 11844
rect 24332 11116 24388 11172
rect 24556 11116 24612 11172
rect 24108 10834 24164 10836
rect 24108 10782 24110 10834
rect 24110 10782 24162 10834
rect 24162 10782 24164 10834
rect 24108 10780 24164 10782
rect 24332 10834 24388 10836
rect 24332 10782 24334 10834
rect 24334 10782 24386 10834
rect 24386 10782 24388 10834
rect 24332 10780 24388 10782
rect 25004 10780 25060 10836
rect 24444 10108 24500 10164
rect 24108 9996 24164 10052
rect 24220 9772 24276 9828
rect 24108 9324 24164 9380
rect 23772 8092 23828 8148
rect 23660 7868 23716 7924
rect 22764 4898 22820 4900
rect 22764 4846 22766 4898
rect 22766 4846 22818 4898
rect 22818 4846 22820 4898
rect 22764 4844 22820 4846
rect 22876 4732 22932 4788
rect 22764 4620 22820 4676
rect 22876 4396 22932 4452
rect 23884 7698 23940 7700
rect 23884 7646 23886 7698
rect 23886 7646 23938 7698
rect 23938 7646 23940 7698
rect 23884 7644 23940 7646
rect 24108 7420 24164 7476
rect 24556 9154 24612 9156
rect 24556 9102 24558 9154
rect 24558 9102 24610 9154
rect 24610 9102 24612 9154
rect 24556 9100 24612 9102
rect 24444 9042 24500 9044
rect 24444 8990 24446 9042
rect 24446 8990 24498 9042
rect 24498 8990 24500 9042
rect 24444 8988 24500 8990
rect 24780 9042 24836 9044
rect 24780 8990 24782 9042
rect 24782 8990 24834 9042
rect 24834 8990 24836 9042
rect 24780 8988 24836 8990
rect 25004 8482 25060 8484
rect 25004 8430 25006 8482
rect 25006 8430 25058 8482
rect 25058 8430 25060 8482
rect 25004 8428 25060 8430
rect 24892 8316 24948 8372
rect 23996 7308 24052 7364
rect 24556 7868 24612 7924
rect 24220 7308 24276 7364
rect 24668 7362 24724 7364
rect 24668 7310 24670 7362
rect 24670 7310 24722 7362
rect 24722 7310 24724 7362
rect 24668 7308 24724 7310
rect 23884 7196 23940 7252
rect 23660 6300 23716 6356
rect 23772 6412 23828 6468
rect 23324 4508 23380 4564
rect 23772 5852 23828 5908
rect 24108 6748 24164 6804
rect 24444 6748 24500 6804
rect 24556 7196 24612 7252
rect 24108 6524 24164 6580
rect 24892 7196 24948 7252
rect 25004 8092 25060 8148
rect 24892 6972 24948 7028
rect 24444 6578 24500 6580
rect 24444 6526 24446 6578
rect 24446 6526 24498 6578
rect 24498 6526 24500 6578
rect 24444 6524 24500 6526
rect 24668 6412 24724 6468
rect 24332 6018 24388 6020
rect 24332 5966 24334 6018
rect 24334 5966 24386 6018
rect 24386 5966 24388 6018
rect 24332 5964 24388 5966
rect 24780 6018 24836 6020
rect 24780 5966 24782 6018
rect 24782 5966 24834 6018
rect 24834 5966 24836 6018
rect 24780 5964 24836 5966
rect 25452 13468 25508 13524
rect 25676 13020 25732 13076
rect 25564 12460 25620 12516
rect 25452 11618 25508 11620
rect 25452 11566 25454 11618
rect 25454 11566 25506 11618
rect 25506 11566 25508 11618
rect 25452 11564 25508 11566
rect 25452 11228 25508 11284
rect 25340 10668 25396 10724
rect 25452 10050 25508 10052
rect 25452 9998 25454 10050
rect 25454 9998 25506 10050
rect 25506 9998 25508 10050
rect 25452 9996 25508 9998
rect 25340 9660 25396 9716
rect 25900 15036 25956 15092
rect 27916 29986 27972 29988
rect 27916 29934 27918 29986
rect 27918 29934 27970 29986
rect 27970 29934 27972 29986
rect 27916 29932 27972 29934
rect 30044 31276 30100 31332
rect 30828 32508 30884 32564
rect 30604 32450 30660 32452
rect 30604 32398 30606 32450
rect 30606 32398 30658 32450
rect 30658 32398 30660 32450
rect 30604 32396 30660 32398
rect 30828 31948 30884 32004
rect 30268 29820 30324 29876
rect 30828 29932 30884 29988
rect 28588 29426 28644 29428
rect 28588 29374 28590 29426
rect 28590 29374 28642 29426
rect 28642 29374 28644 29426
rect 28588 29372 28644 29374
rect 29148 29372 29204 29428
rect 29484 28642 29540 28644
rect 29484 28590 29486 28642
rect 29486 28590 29538 28642
rect 29538 28590 29540 28642
rect 29484 28588 29540 28590
rect 28588 28028 28644 28084
rect 31836 31276 31892 31332
rect 31948 31052 32004 31108
rect 31836 30156 31892 30212
rect 32060 30156 32116 30212
rect 31612 29650 31668 29652
rect 31612 29598 31614 29650
rect 31614 29598 31666 29650
rect 31666 29598 31668 29650
rect 31612 29596 31668 29598
rect 31052 28642 31108 28644
rect 31052 28590 31054 28642
rect 31054 28590 31106 28642
rect 31106 28590 31108 28642
rect 31052 28588 31108 28590
rect 32172 29596 32228 29652
rect 31948 28700 32004 28756
rect 29036 28082 29092 28084
rect 29036 28030 29038 28082
rect 29038 28030 29090 28082
rect 29090 28030 29092 28082
rect 29036 28028 29092 28030
rect 27804 27692 27860 27748
rect 27804 27020 27860 27076
rect 27580 25340 27636 25396
rect 27692 25228 27748 25284
rect 28252 27692 28308 27748
rect 28476 27468 28532 27524
rect 28924 27580 28980 27636
rect 27916 25900 27972 25956
rect 28588 26796 28644 26852
rect 27916 25340 27972 25396
rect 27468 23212 27524 23268
rect 27580 23100 27636 23156
rect 26908 21868 26964 21924
rect 26796 21420 26852 21476
rect 27244 21474 27300 21476
rect 27244 21422 27246 21474
rect 27246 21422 27298 21474
rect 27298 21422 27300 21474
rect 27244 21420 27300 21422
rect 26796 20412 26852 20468
rect 26236 20076 26292 20132
rect 26236 19740 26292 19796
rect 26236 19234 26292 19236
rect 26236 19182 26238 19234
rect 26238 19182 26290 19234
rect 26290 19182 26292 19234
rect 26236 19180 26292 19182
rect 26236 17724 26292 17780
rect 26236 17164 26292 17220
rect 26236 16940 26292 16996
rect 26460 19516 26516 19572
rect 26684 19516 26740 19572
rect 27244 20636 27300 20692
rect 27132 19292 27188 19348
rect 26908 17666 26964 17668
rect 26908 17614 26910 17666
rect 26910 17614 26962 17666
rect 26962 17614 26964 17666
rect 26908 17612 26964 17614
rect 26572 17500 26628 17556
rect 26908 17388 26964 17444
rect 26572 15314 26628 15316
rect 26572 15262 26574 15314
rect 26574 15262 26626 15314
rect 26626 15262 26628 15314
rect 26572 15260 26628 15262
rect 26796 16658 26852 16660
rect 26796 16606 26798 16658
rect 26798 16606 26850 16658
rect 26850 16606 26852 16658
rect 26796 16604 26852 16606
rect 26684 16044 26740 16100
rect 26460 15148 26516 15204
rect 26236 14418 26292 14420
rect 26236 14366 26238 14418
rect 26238 14366 26290 14418
rect 26290 14366 26292 14418
rect 26236 14364 26292 14366
rect 25788 11788 25844 11844
rect 26124 12290 26180 12292
rect 26124 12238 26126 12290
rect 26126 12238 26178 12290
rect 26178 12238 26180 12290
rect 26124 12236 26180 12238
rect 25900 11564 25956 11620
rect 25676 11506 25732 11508
rect 25676 11454 25678 11506
rect 25678 11454 25730 11506
rect 25730 11454 25732 11506
rect 25676 11452 25732 11454
rect 25788 11170 25844 11172
rect 25788 11118 25790 11170
rect 25790 11118 25842 11170
rect 25842 11118 25844 11170
rect 25788 11116 25844 11118
rect 25788 10722 25844 10724
rect 25788 10670 25790 10722
rect 25790 10670 25842 10722
rect 25842 10670 25844 10722
rect 25788 10668 25844 10670
rect 25676 10556 25732 10612
rect 26012 10556 26068 10612
rect 26348 13580 26404 13636
rect 26572 14140 26628 14196
rect 26796 16268 26852 16324
rect 27132 18732 27188 18788
rect 27244 17052 27300 17108
rect 27132 16882 27188 16884
rect 27132 16830 27134 16882
rect 27134 16830 27186 16882
rect 27186 16830 27188 16882
rect 27132 16828 27188 16830
rect 26908 15426 26964 15428
rect 26908 15374 26910 15426
rect 26910 15374 26962 15426
rect 26962 15374 26964 15426
rect 26908 15372 26964 15374
rect 26908 14588 26964 14644
rect 27132 15820 27188 15876
rect 27132 14418 27188 14420
rect 27132 14366 27134 14418
rect 27134 14366 27186 14418
rect 27186 14366 27188 14418
rect 27132 14364 27188 14366
rect 26908 13244 26964 13300
rect 26572 11788 26628 11844
rect 26572 11340 26628 11396
rect 25340 8652 25396 8708
rect 25228 8316 25284 8372
rect 25340 7586 25396 7588
rect 25340 7534 25342 7586
rect 25342 7534 25394 7586
rect 25394 7534 25396 7586
rect 25340 7532 25396 7534
rect 25340 6972 25396 7028
rect 25340 6188 25396 6244
rect 25788 9324 25844 9380
rect 25676 9042 25732 9044
rect 25676 8990 25678 9042
rect 25678 8990 25730 9042
rect 25730 8990 25732 9042
rect 25676 8988 25732 8990
rect 25788 8540 25844 8596
rect 26572 9660 26628 9716
rect 26460 9324 26516 9380
rect 26124 9212 26180 9268
rect 26572 9154 26628 9156
rect 26572 9102 26574 9154
rect 26574 9102 26626 9154
rect 26626 9102 26628 9154
rect 26572 9100 26628 9102
rect 26012 8652 26068 8708
rect 25788 8092 25844 8148
rect 26348 8034 26404 8036
rect 26348 7982 26350 8034
rect 26350 7982 26402 8034
rect 26402 7982 26404 8034
rect 26348 7980 26404 7982
rect 26012 7586 26068 7588
rect 26012 7534 26014 7586
rect 26014 7534 26066 7586
rect 26066 7534 26068 7586
rect 26012 7532 26068 7534
rect 26236 7474 26292 7476
rect 26236 7422 26238 7474
rect 26238 7422 26290 7474
rect 26290 7422 26292 7474
rect 26236 7420 26292 7422
rect 26012 7362 26068 7364
rect 26012 7310 26014 7362
rect 26014 7310 26066 7362
rect 26066 7310 26068 7362
rect 26012 7308 26068 7310
rect 25676 6972 25732 7028
rect 25900 7084 25956 7140
rect 24108 5404 24164 5460
rect 24780 5516 24836 5572
rect 24332 5292 24388 5348
rect 24332 4562 24388 4564
rect 24332 4510 24334 4562
rect 24334 4510 24386 4562
rect 24386 4510 24388 4562
rect 24332 4508 24388 4510
rect 23100 4060 23156 4116
rect 21980 3554 22036 3556
rect 21980 3502 21982 3554
rect 21982 3502 22034 3554
rect 22034 3502 22036 3554
rect 21980 3500 22036 3502
rect 23100 3500 23156 3556
rect 19740 3276 19796 3332
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 25228 5292 25284 5348
rect 25452 5292 25508 5348
rect 25116 5068 25172 5124
rect 25452 4956 25508 5012
rect 25340 4620 25396 4676
rect 25452 4562 25508 4564
rect 25452 4510 25454 4562
rect 25454 4510 25506 4562
rect 25506 4510 25508 4562
rect 25452 4508 25508 4510
rect 25228 4450 25284 4452
rect 25228 4398 25230 4450
rect 25230 4398 25282 4450
rect 25282 4398 25284 4450
rect 25228 4396 25284 4398
rect 25788 6300 25844 6356
rect 26908 11900 26964 11956
rect 27020 11004 27076 11060
rect 27244 13132 27300 13188
rect 28140 25900 28196 25956
rect 28476 26066 28532 26068
rect 28476 26014 28478 26066
rect 28478 26014 28530 26066
rect 28530 26014 28532 26066
rect 28476 26012 28532 26014
rect 28252 25452 28308 25508
rect 29148 27074 29204 27076
rect 29148 27022 29150 27074
rect 29150 27022 29202 27074
rect 29202 27022 29204 27074
rect 29148 27020 29204 27022
rect 29820 28082 29876 28084
rect 29820 28030 29822 28082
rect 29822 28030 29874 28082
rect 29874 28030 29876 28082
rect 29820 28028 29876 28030
rect 29260 26962 29316 26964
rect 29260 26910 29262 26962
rect 29262 26910 29314 26962
rect 29314 26910 29316 26962
rect 29260 26908 29316 26910
rect 29148 25788 29204 25844
rect 30940 28028 30996 28084
rect 31276 28364 31332 28420
rect 34076 35138 34132 35140
rect 34076 35086 34078 35138
rect 34078 35086 34130 35138
rect 34130 35086 34132 35138
rect 34076 35084 34132 35086
rect 33516 34972 33572 35028
rect 32732 34802 32788 34804
rect 32732 34750 32734 34802
rect 32734 34750 32786 34802
rect 32786 34750 32788 34802
rect 32732 34748 32788 34750
rect 34860 36652 34916 36708
rect 34860 35922 34916 35924
rect 34860 35870 34862 35922
rect 34862 35870 34914 35922
rect 34914 35870 34916 35922
rect 34860 35868 34916 35870
rect 34300 35474 34356 35476
rect 34300 35422 34302 35474
rect 34302 35422 34354 35474
rect 34354 35422 34356 35474
rect 34300 35420 34356 35422
rect 34524 35698 34580 35700
rect 34524 35646 34526 35698
rect 34526 35646 34578 35698
rect 34578 35646 34580 35698
rect 34524 35644 34580 35646
rect 34412 35308 34468 35364
rect 34076 34524 34132 34580
rect 33516 34300 33572 34356
rect 34188 34354 34244 34356
rect 34188 34302 34190 34354
rect 34190 34302 34242 34354
rect 34242 34302 34244 34354
rect 34188 34300 34244 34302
rect 33628 34242 33684 34244
rect 33628 34190 33630 34242
rect 33630 34190 33682 34242
rect 33682 34190 33684 34242
rect 33628 34188 33684 34190
rect 32844 34076 32900 34132
rect 34412 34076 34468 34132
rect 35644 38668 35700 38724
rect 35756 37772 35812 37828
rect 35532 37548 35588 37604
rect 35644 37436 35700 37492
rect 35084 37324 35140 37380
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35420 36706 35476 36708
rect 35420 36654 35422 36706
rect 35422 36654 35474 36706
rect 35474 36654 35476 36706
rect 35420 36652 35476 36654
rect 35196 36092 35252 36148
rect 36092 37884 36148 37940
rect 35980 37660 36036 37716
rect 36092 36706 36148 36708
rect 36092 36654 36094 36706
rect 36094 36654 36146 36706
rect 36146 36654 36148 36706
rect 36092 36652 36148 36654
rect 35980 36370 36036 36372
rect 35980 36318 35982 36370
rect 35982 36318 36034 36370
rect 36034 36318 36036 36370
rect 35980 36316 36036 36318
rect 35868 35756 35924 35812
rect 36092 35644 36148 35700
rect 36204 35868 36260 35924
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35756 35308 35812 35364
rect 34972 34300 35028 34356
rect 34860 34242 34916 34244
rect 34860 34190 34862 34242
rect 34862 34190 34914 34242
rect 34914 34190 34916 34242
rect 34860 34188 34916 34190
rect 34748 34130 34804 34132
rect 34748 34078 34750 34130
rect 34750 34078 34802 34130
rect 34802 34078 34804 34130
rect 34748 34076 34804 34078
rect 36316 34860 36372 34916
rect 36428 33852 36484 33908
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 34300 33292 34356 33348
rect 36204 32732 36260 32788
rect 32732 31948 32788 32004
rect 32956 31612 33012 31668
rect 32956 31052 33012 31108
rect 32396 28252 32452 28308
rect 32620 30156 32676 30212
rect 32732 30044 32788 30100
rect 33180 31276 33236 31332
rect 33068 29372 33124 29428
rect 33740 31612 33796 31668
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 34188 31778 34244 31780
rect 34188 31726 34190 31778
rect 34190 31726 34242 31778
rect 34242 31726 34244 31778
rect 34188 31724 34244 31726
rect 33628 31276 33684 31332
rect 37100 44380 37156 44436
rect 37884 48914 37940 48916
rect 37884 48862 37886 48914
rect 37886 48862 37938 48914
rect 37938 48862 37940 48914
rect 37884 48860 37940 48862
rect 38444 49084 38500 49140
rect 38332 48914 38388 48916
rect 38332 48862 38334 48914
rect 38334 48862 38386 48914
rect 38386 48862 38388 48914
rect 38332 48860 38388 48862
rect 38220 48412 38276 48468
rect 37436 47458 37492 47460
rect 37436 47406 37438 47458
rect 37438 47406 37490 47458
rect 37490 47406 37492 47458
rect 37436 47404 37492 47406
rect 37660 48130 37716 48132
rect 37660 48078 37662 48130
rect 37662 48078 37714 48130
rect 37714 48078 37716 48130
rect 37660 48076 37716 48078
rect 38556 48412 38612 48468
rect 38108 47964 38164 48020
rect 38668 48018 38724 48020
rect 38668 47966 38670 48018
rect 38670 47966 38722 48018
rect 38722 47966 38724 48018
rect 38668 47964 38724 47966
rect 38220 47404 38276 47460
rect 38444 46956 38500 47012
rect 37996 46562 38052 46564
rect 37996 46510 37998 46562
rect 37998 46510 38050 46562
rect 38050 46510 38052 46562
rect 37996 46508 38052 46510
rect 38444 46562 38500 46564
rect 38444 46510 38446 46562
rect 38446 46510 38498 46562
rect 38498 46510 38500 46562
rect 38444 46508 38500 46510
rect 37548 44156 37604 44212
rect 37436 43596 37492 43652
rect 36988 40572 37044 40628
rect 37548 43484 37604 43540
rect 37212 40908 37268 40964
rect 38780 46956 38836 47012
rect 38780 45666 38836 45668
rect 38780 45614 38782 45666
rect 38782 45614 38834 45666
rect 38834 45614 38836 45666
rect 38780 45612 38836 45614
rect 39004 48466 39060 48468
rect 39004 48414 39006 48466
rect 39006 48414 39058 48466
rect 39058 48414 39060 48466
rect 39004 48412 39060 48414
rect 40236 49810 40292 49812
rect 40236 49758 40238 49810
rect 40238 49758 40290 49810
rect 40290 49758 40292 49810
rect 40236 49756 40292 49758
rect 40460 50204 40516 50260
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 45724 56252 45780 56308
rect 48412 56306 48468 56308
rect 48412 56254 48414 56306
rect 48414 56254 48466 56306
rect 48466 56254 48468 56306
rect 48412 56252 48468 56254
rect 41692 56028 41748 56084
rect 42588 56082 42644 56084
rect 42588 56030 42590 56082
rect 42590 56030 42642 56082
rect 42642 56030 42644 56082
rect 42588 56028 42644 56030
rect 46508 56028 46564 56084
rect 41804 55244 41860 55300
rect 40684 53954 40740 53956
rect 40684 53902 40686 53954
rect 40686 53902 40738 53954
rect 40738 53902 40740 53954
rect 40684 53900 40740 53902
rect 43372 55298 43428 55300
rect 43372 55246 43374 55298
rect 43374 55246 43426 55298
rect 43426 55246 43428 55298
rect 43372 55244 43428 55246
rect 42476 55186 42532 55188
rect 42476 55134 42478 55186
rect 42478 55134 42530 55186
rect 42530 55134 42532 55186
rect 42476 55132 42532 55134
rect 42700 55186 42756 55188
rect 42700 55134 42702 55186
rect 42702 55134 42754 55186
rect 42754 55134 42756 55186
rect 42700 55132 42756 55134
rect 43820 55132 43876 55188
rect 42588 55074 42644 55076
rect 42588 55022 42590 55074
rect 42590 55022 42642 55074
rect 42642 55022 42644 55074
rect 42588 55020 42644 55022
rect 41916 54236 41972 54292
rect 42140 54514 42196 54516
rect 42140 54462 42142 54514
rect 42142 54462 42194 54514
rect 42194 54462 42196 54514
rect 42140 54460 42196 54462
rect 42700 54348 42756 54404
rect 42812 54460 42868 54516
rect 42028 53900 42084 53956
rect 43708 54514 43764 54516
rect 43708 54462 43710 54514
rect 43710 54462 43762 54514
rect 43762 54462 43764 54514
rect 43708 54460 43764 54462
rect 40796 53842 40852 53844
rect 40796 53790 40798 53842
rect 40798 53790 40850 53842
rect 40850 53790 40852 53842
rect 40796 53788 40852 53790
rect 42252 53730 42308 53732
rect 42252 53678 42254 53730
rect 42254 53678 42306 53730
rect 42306 53678 42308 53730
rect 42252 53676 42308 53678
rect 41356 53618 41412 53620
rect 41356 53566 41358 53618
rect 41358 53566 41410 53618
rect 41410 53566 41412 53618
rect 41356 53564 41412 53566
rect 43260 53676 43316 53732
rect 42476 53564 42532 53620
rect 41244 52332 41300 52388
rect 41020 52220 41076 52276
rect 41132 52162 41188 52164
rect 41132 52110 41134 52162
rect 41134 52110 41186 52162
rect 41186 52110 41188 52162
rect 41132 52108 41188 52110
rect 41692 52386 41748 52388
rect 41692 52334 41694 52386
rect 41694 52334 41746 52386
rect 41746 52334 41748 52386
rect 41692 52332 41748 52334
rect 40908 51548 40964 51604
rect 41692 51212 41748 51268
rect 40572 49980 40628 50036
rect 41020 50204 41076 50260
rect 41468 50034 41524 50036
rect 41468 49982 41470 50034
rect 41470 49982 41522 50034
rect 41522 49982 41524 50034
rect 41468 49980 41524 49982
rect 40348 49196 40404 49252
rect 39564 49026 39620 49028
rect 39564 48974 39566 49026
rect 39566 48974 39618 49026
rect 39618 48974 39620 49026
rect 39564 48972 39620 48974
rect 39900 48914 39956 48916
rect 39900 48862 39902 48914
rect 39902 48862 39954 48914
rect 39954 48862 39956 48914
rect 39900 48860 39956 48862
rect 40908 48972 40964 49028
rect 40460 48802 40516 48804
rect 40460 48750 40462 48802
rect 40462 48750 40514 48802
rect 40514 48750 40516 48802
rect 40460 48748 40516 48750
rect 39452 48130 39508 48132
rect 39452 48078 39454 48130
rect 39454 48078 39506 48130
rect 39506 48078 39508 48130
rect 39452 48076 39508 48078
rect 39340 47570 39396 47572
rect 39340 47518 39342 47570
rect 39342 47518 39394 47570
rect 39394 47518 39396 47570
rect 39340 47516 39396 47518
rect 40348 47964 40404 48020
rect 40236 47516 40292 47572
rect 37772 43538 37828 43540
rect 37772 43486 37774 43538
rect 37774 43486 37826 43538
rect 37826 43486 37828 43538
rect 37772 43484 37828 43486
rect 38220 44434 38276 44436
rect 38220 44382 38222 44434
rect 38222 44382 38274 44434
rect 38274 44382 38276 44434
rect 38220 44380 38276 44382
rect 37996 44268 38052 44324
rect 38332 44268 38388 44324
rect 39004 44322 39060 44324
rect 39004 44270 39006 44322
rect 39006 44270 39058 44322
rect 39058 44270 39060 44322
rect 39004 44268 39060 44270
rect 38668 43596 38724 43652
rect 37996 42812 38052 42868
rect 38556 43426 38612 43428
rect 38556 43374 38558 43426
rect 38558 43374 38610 43426
rect 38610 43374 38612 43426
rect 38556 43372 38612 43374
rect 37884 42642 37940 42644
rect 37884 42590 37886 42642
rect 37886 42590 37938 42642
rect 37938 42590 37940 42642
rect 37884 42588 37940 42590
rect 38556 42476 38612 42532
rect 38892 42476 38948 42532
rect 37996 41804 38052 41860
rect 38668 41020 38724 41076
rect 36988 37436 37044 37492
rect 36764 35922 36820 35924
rect 36764 35870 36766 35922
rect 36766 35870 36818 35922
rect 36818 35870 36820 35922
rect 36764 35868 36820 35870
rect 36652 35084 36708 35140
rect 37548 37884 37604 37940
rect 37660 37490 37716 37492
rect 37660 37438 37662 37490
rect 37662 37438 37714 37490
rect 37714 37438 37716 37490
rect 37660 37436 37716 37438
rect 38780 40348 38836 40404
rect 38332 38722 38388 38724
rect 38332 38670 38334 38722
rect 38334 38670 38386 38722
rect 38386 38670 38388 38722
rect 38332 38668 38388 38670
rect 37884 37826 37940 37828
rect 37884 37774 37886 37826
rect 37886 37774 37938 37826
rect 37938 37774 37940 37826
rect 37884 37772 37940 37774
rect 38108 37324 38164 37380
rect 38444 37378 38500 37380
rect 38444 37326 38446 37378
rect 38446 37326 38498 37378
rect 38498 37326 38500 37378
rect 38444 37324 38500 37326
rect 37436 35810 37492 35812
rect 37436 35758 37438 35810
rect 37438 35758 37490 35810
rect 37490 35758 37492 35810
rect 37436 35756 37492 35758
rect 37548 35698 37604 35700
rect 37548 35646 37550 35698
rect 37550 35646 37602 35698
rect 37602 35646 37604 35698
rect 37548 35644 37604 35646
rect 37996 35308 38052 35364
rect 38108 35756 38164 35812
rect 37324 35196 37380 35252
rect 37324 34914 37380 34916
rect 37324 34862 37326 34914
rect 37326 34862 37378 34914
rect 37378 34862 37380 34914
rect 37324 34860 37380 34862
rect 38220 33852 38276 33908
rect 38220 33404 38276 33460
rect 37548 32956 37604 33012
rect 37212 32786 37268 32788
rect 37212 32734 37214 32786
rect 37214 32734 37266 32786
rect 37266 32734 37268 32786
rect 37212 32732 37268 32734
rect 36652 32620 36708 32676
rect 37324 32620 37380 32676
rect 37212 32508 37268 32564
rect 36540 31164 36596 31220
rect 33628 31052 33684 31108
rect 33964 31052 34020 31108
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 33964 30210 34020 30212
rect 33964 30158 33966 30210
rect 33966 30158 34018 30210
rect 34018 30158 34020 30210
rect 33964 30156 34020 30158
rect 33292 30098 33348 30100
rect 33292 30046 33294 30098
rect 33294 30046 33346 30098
rect 33346 30046 33348 30098
rect 33292 30044 33348 30046
rect 33404 29596 33460 29652
rect 33292 28812 33348 28868
rect 33180 28700 33236 28756
rect 37772 32674 37828 32676
rect 37772 32622 37774 32674
rect 37774 32622 37826 32674
rect 37826 32622 37828 32674
rect 37772 32620 37828 32622
rect 38108 32732 38164 32788
rect 38780 35698 38836 35700
rect 38780 35646 38782 35698
rect 38782 35646 38834 35698
rect 38834 35646 38836 35698
rect 38780 35644 38836 35646
rect 38668 35308 38724 35364
rect 38556 34802 38612 34804
rect 38556 34750 38558 34802
rect 38558 34750 38610 34802
rect 38610 34750 38612 34802
rect 38556 34748 38612 34750
rect 39228 45778 39284 45780
rect 39228 45726 39230 45778
rect 39230 45726 39282 45778
rect 39282 45726 39284 45778
rect 39228 45724 39284 45726
rect 39340 45388 39396 45444
rect 40124 46898 40180 46900
rect 40124 46846 40126 46898
rect 40126 46846 40178 46898
rect 40178 46846 40180 46898
rect 40124 46844 40180 46846
rect 39900 46620 39956 46676
rect 40012 45724 40068 45780
rect 39676 43484 39732 43540
rect 39788 45612 39844 45668
rect 39340 43260 39396 43316
rect 40796 47964 40852 48020
rect 43148 53618 43204 53620
rect 43148 53566 43150 53618
rect 43150 53566 43202 53618
rect 43202 53566 43204 53618
rect 43148 53564 43204 53566
rect 42476 52332 42532 52388
rect 44492 54402 44548 54404
rect 44492 54350 44494 54402
rect 44494 54350 44546 54402
rect 44546 54350 44548 54402
rect 44492 54348 44548 54350
rect 47404 56082 47460 56084
rect 47404 56030 47406 56082
rect 47406 56030 47458 56082
rect 47458 56030 47460 56082
rect 47404 56028 47460 56030
rect 53004 56028 53060 56084
rect 45500 54738 45556 54740
rect 45500 54686 45502 54738
rect 45502 54686 45554 54738
rect 45554 54686 45556 54738
rect 45500 54684 45556 54686
rect 46396 54572 46452 54628
rect 46956 54626 47012 54628
rect 46956 54574 46958 54626
rect 46958 54574 47010 54626
rect 47010 54574 47012 54626
rect 46956 54572 47012 54574
rect 44940 54236 44996 54292
rect 46844 53900 46900 53956
rect 46508 53788 46564 53844
rect 45836 53676 45892 53732
rect 43932 52332 43988 52388
rect 43260 52274 43316 52276
rect 43260 52222 43262 52274
rect 43262 52222 43314 52274
rect 43314 52222 43316 52274
rect 43260 52220 43316 52222
rect 43484 52220 43540 52276
rect 43260 51996 43316 52052
rect 42700 51884 42756 51940
rect 42476 51660 42532 51716
rect 43036 51100 43092 51156
rect 44044 52274 44100 52276
rect 44044 52222 44046 52274
rect 44046 52222 44098 52274
rect 44098 52222 44100 52274
rect 44044 52220 44100 52222
rect 45164 52220 45220 52276
rect 43596 52162 43652 52164
rect 43596 52110 43598 52162
rect 43598 52110 43650 52162
rect 43650 52110 43652 52162
rect 43596 52108 43652 52110
rect 43484 52050 43540 52052
rect 43484 51998 43486 52050
rect 43486 51998 43538 52050
rect 43538 51998 43540 52050
rect 43484 51996 43540 51998
rect 42700 50988 42756 51044
rect 42140 50204 42196 50260
rect 43484 50988 43540 51044
rect 43260 50540 43316 50596
rect 42812 50370 42868 50372
rect 42812 50318 42814 50370
rect 42814 50318 42866 50370
rect 42866 50318 42868 50370
rect 42812 50316 42868 50318
rect 43372 50204 43428 50260
rect 43372 49868 43428 49924
rect 44828 52162 44884 52164
rect 44828 52110 44830 52162
rect 44830 52110 44882 52162
rect 44882 52110 44884 52162
rect 44828 52108 44884 52110
rect 45612 52444 45668 52500
rect 43708 51154 43764 51156
rect 43708 51102 43710 51154
rect 43710 51102 43762 51154
rect 43762 51102 43764 51154
rect 43708 51100 43764 51102
rect 43596 50316 43652 50372
rect 47068 53788 47124 53844
rect 47180 53730 47236 53732
rect 47180 53678 47182 53730
rect 47182 53678 47234 53730
rect 47234 53678 47236 53730
rect 47180 53676 47236 53678
rect 46172 52332 46228 52388
rect 48188 55020 48244 55076
rect 48748 55020 48804 55076
rect 47628 54514 47684 54516
rect 47628 54462 47630 54514
rect 47630 54462 47682 54514
rect 47682 54462 47684 54514
rect 47628 54460 47684 54462
rect 47516 53900 47572 53956
rect 47852 54290 47908 54292
rect 47852 54238 47854 54290
rect 47854 54238 47906 54290
rect 47906 54238 47908 54290
rect 47852 54236 47908 54238
rect 47740 53788 47796 53844
rect 48300 54514 48356 54516
rect 48300 54462 48302 54514
rect 48302 54462 48354 54514
rect 48354 54462 48356 54514
rect 48300 54460 48356 54462
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 50764 54684 50820 54740
rect 49084 54626 49140 54628
rect 49084 54574 49086 54626
rect 49086 54574 49138 54626
rect 49138 54574 49140 54626
rect 49084 54572 49140 54574
rect 48972 54514 49028 54516
rect 48972 54462 48974 54514
rect 48974 54462 49026 54514
rect 49026 54462 49028 54514
rect 48972 54460 49028 54462
rect 49532 54514 49588 54516
rect 49532 54462 49534 54514
rect 49534 54462 49586 54514
rect 49586 54462 49588 54514
rect 49532 54460 49588 54462
rect 49196 54348 49252 54404
rect 48076 53900 48132 53956
rect 47628 53618 47684 53620
rect 47628 53566 47630 53618
rect 47630 53566 47682 53618
rect 47682 53566 47684 53618
rect 47628 53564 47684 53566
rect 47404 52220 47460 52276
rect 45836 51212 45892 51268
rect 46508 51266 46564 51268
rect 46508 51214 46510 51266
rect 46510 51214 46562 51266
rect 46562 51214 46564 51266
rect 46508 51212 46564 51214
rect 47068 51548 47124 51604
rect 46956 51266 47012 51268
rect 46956 51214 46958 51266
rect 46958 51214 47010 51266
rect 47010 51214 47012 51266
rect 46956 51212 47012 51214
rect 45612 50594 45668 50596
rect 45612 50542 45614 50594
rect 45614 50542 45666 50594
rect 45666 50542 45668 50594
rect 45612 50540 45668 50542
rect 44268 50482 44324 50484
rect 44268 50430 44270 50482
rect 44270 50430 44322 50482
rect 44322 50430 44324 50482
rect 44268 50428 44324 50430
rect 44380 49980 44436 50036
rect 43820 49026 43876 49028
rect 43820 48974 43822 49026
rect 43822 48974 43874 49026
rect 43874 48974 43876 49026
rect 43820 48972 43876 48974
rect 44268 49196 44324 49252
rect 43596 48914 43652 48916
rect 43596 48862 43598 48914
rect 43598 48862 43650 48914
rect 43650 48862 43652 48914
rect 43596 48860 43652 48862
rect 40908 46674 40964 46676
rect 40908 46622 40910 46674
rect 40910 46622 40962 46674
rect 40962 46622 40964 46674
rect 40908 46620 40964 46622
rect 41244 46620 41300 46676
rect 41580 46844 41636 46900
rect 41244 46114 41300 46116
rect 41244 46062 41246 46114
rect 41246 46062 41298 46114
rect 41298 46062 41300 46114
rect 41244 46060 41300 46062
rect 40124 44716 40180 44772
rect 40348 43484 40404 43540
rect 40236 41916 40292 41972
rect 39676 41186 39732 41188
rect 39676 41134 39678 41186
rect 39678 41134 39730 41186
rect 39730 41134 39732 41186
rect 39676 41132 39732 41134
rect 39900 39394 39956 39396
rect 39900 39342 39902 39394
rect 39902 39342 39954 39394
rect 39954 39342 39956 39394
rect 39900 39340 39956 39342
rect 39228 38722 39284 38724
rect 39228 38670 39230 38722
rect 39230 38670 39282 38722
rect 39282 38670 39284 38722
rect 39228 38668 39284 38670
rect 39004 37772 39060 37828
rect 39116 37436 39172 37492
rect 39788 37436 39844 37492
rect 39340 37378 39396 37380
rect 39340 37326 39342 37378
rect 39342 37326 39394 37378
rect 39394 37326 39396 37378
rect 39340 37324 39396 37326
rect 41020 44716 41076 44772
rect 41356 44492 41412 44548
rect 41916 46956 41972 47012
rect 42252 46620 42308 46676
rect 41916 45724 41972 45780
rect 42140 46060 42196 46116
rect 41468 44044 41524 44100
rect 40908 43538 40964 43540
rect 40908 43486 40910 43538
rect 40910 43486 40962 43538
rect 40962 43486 40964 43538
rect 40908 43484 40964 43486
rect 41804 43484 41860 43540
rect 42028 44044 42084 44100
rect 41916 42588 41972 42644
rect 42924 46674 42980 46676
rect 42924 46622 42926 46674
rect 42926 46622 42978 46674
rect 42978 46622 42980 46674
rect 42924 46620 42980 46622
rect 42476 45388 42532 45444
rect 43372 45164 43428 45220
rect 43484 44828 43540 44884
rect 42700 44322 42756 44324
rect 42700 44270 42702 44322
rect 42702 44270 42754 44322
rect 42754 44270 42756 44322
rect 42700 44268 42756 44270
rect 43484 44098 43540 44100
rect 43484 44046 43486 44098
rect 43486 44046 43538 44098
rect 43538 44046 43540 44098
rect 43484 44044 43540 44046
rect 42588 43538 42644 43540
rect 42588 43486 42590 43538
rect 42590 43486 42642 43538
rect 42642 43486 42644 43538
rect 42588 43484 42644 43486
rect 42924 43484 42980 43540
rect 42028 41916 42084 41972
rect 39228 33516 39284 33572
rect 38668 33404 38724 33460
rect 37548 32562 37604 32564
rect 37548 32510 37550 32562
rect 37550 32510 37602 32562
rect 37602 32510 37604 32562
rect 37548 32508 37604 32510
rect 38332 31164 38388 31220
rect 36316 29650 36372 29652
rect 36316 29598 36318 29650
rect 36318 29598 36370 29650
rect 36370 29598 36372 29650
rect 36316 29596 36372 29598
rect 38668 31778 38724 31780
rect 38668 31726 38670 31778
rect 38670 31726 38722 31778
rect 38722 31726 38724 31778
rect 38668 31724 38724 31726
rect 38780 31218 38836 31220
rect 38780 31166 38782 31218
rect 38782 31166 38834 31218
rect 38834 31166 38836 31218
rect 38780 31164 38836 31166
rect 39564 36258 39620 36260
rect 39564 36206 39566 36258
rect 39566 36206 39618 36258
rect 39618 36206 39620 36258
rect 39564 36204 39620 36206
rect 41692 41186 41748 41188
rect 41692 41134 41694 41186
rect 41694 41134 41746 41186
rect 41746 41134 41748 41186
rect 41692 41132 41748 41134
rect 41804 40626 41860 40628
rect 41804 40574 41806 40626
rect 41806 40574 41858 40626
rect 41858 40574 41860 40626
rect 41804 40572 41860 40574
rect 42028 41410 42084 41412
rect 42028 41358 42030 41410
rect 42030 41358 42082 41410
rect 42082 41358 42084 41410
rect 42028 41356 42084 41358
rect 42588 42642 42644 42644
rect 42588 42590 42590 42642
rect 42590 42590 42642 42642
rect 42642 42590 42644 42642
rect 42588 42588 42644 42590
rect 42476 41970 42532 41972
rect 42476 41918 42478 41970
rect 42478 41918 42530 41970
rect 42530 41918 42532 41970
rect 42476 41916 42532 41918
rect 41580 39116 41636 39172
rect 41804 39340 41860 39396
rect 41580 38780 41636 38836
rect 41580 38220 41636 38276
rect 41356 37884 41412 37940
rect 41020 37660 41076 37716
rect 42364 39116 42420 39172
rect 42140 38834 42196 38836
rect 42140 38782 42142 38834
rect 42142 38782 42194 38834
rect 42194 38782 42196 38834
rect 42140 38780 42196 38782
rect 42252 37938 42308 37940
rect 42252 37886 42254 37938
rect 42254 37886 42306 37938
rect 42306 37886 42308 37938
rect 42252 37884 42308 37886
rect 41020 36988 41076 37044
rect 40908 36204 40964 36260
rect 41244 36540 41300 36596
rect 42700 39394 42756 39396
rect 42700 39342 42702 39394
rect 42702 39342 42754 39394
rect 42754 39342 42756 39394
rect 42700 39340 42756 39342
rect 42588 38892 42644 38948
rect 43484 43372 43540 43428
rect 42924 42588 42980 42644
rect 43596 42588 43652 42644
rect 43036 39116 43092 39172
rect 43260 38834 43316 38836
rect 43260 38782 43262 38834
rect 43262 38782 43314 38834
rect 43314 38782 43316 38834
rect 43260 38780 43316 38782
rect 42812 37996 42868 38052
rect 42028 37042 42084 37044
rect 42028 36990 42030 37042
rect 42030 36990 42082 37042
rect 42082 36990 42084 37042
rect 42028 36988 42084 36990
rect 41804 36594 41860 36596
rect 41804 36542 41806 36594
rect 41806 36542 41858 36594
rect 41858 36542 41860 36594
rect 41804 36540 41860 36542
rect 42364 36204 42420 36260
rect 39452 35644 39508 35700
rect 43036 36204 43092 36260
rect 40572 35026 40628 35028
rect 40572 34974 40574 35026
rect 40574 34974 40626 35026
rect 40626 34974 40628 35026
rect 40572 34972 40628 34974
rect 39788 33516 39844 33572
rect 39004 31218 39060 31220
rect 39004 31166 39006 31218
rect 39006 31166 39058 31218
rect 39058 31166 39060 31218
rect 39004 31164 39060 31166
rect 40908 33516 40964 33572
rect 40460 33404 40516 33460
rect 38892 30434 38948 30436
rect 38892 30382 38894 30434
rect 38894 30382 38946 30434
rect 38946 30382 38948 30434
rect 38892 30380 38948 30382
rect 41020 32172 41076 32228
rect 43260 38050 43316 38052
rect 43260 37998 43262 38050
rect 43262 37998 43314 38050
rect 43314 37998 43316 38050
rect 43260 37996 43316 37998
rect 43596 39058 43652 39060
rect 43596 39006 43598 39058
rect 43598 39006 43650 39058
rect 43650 39006 43652 39058
rect 43596 39004 43652 39006
rect 45276 49868 45332 49924
rect 44940 48188 44996 48244
rect 44044 47068 44100 47124
rect 44156 46956 44212 47012
rect 45164 46844 45220 46900
rect 45388 49084 45444 49140
rect 45612 48972 45668 49028
rect 45612 48188 45668 48244
rect 45164 45218 45220 45220
rect 45164 45166 45166 45218
rect 45166 45166 45218 45218
rect 45218 45166 45220 45218
rect 45164 45164 45220 45166
rect 44940 44828 44996 44884
rect 45388 45052 45444 45108
rect 45276 44828 45332 44884
rect 44828 44098 44884 44100
rect 44828 44046 44830 44098
rect 44830 44046 44882 44098
rect 44882 44046 44884 44098
rect 44828 44044 44884 44046
rect 44380 43538 44436 43540
rect 44380 43486 44382 43538
rect 44382 43486 44434 43538
rect 44434 43486 44436 43538
rect 44380 43484 44436 43486
rect 45276 44268 45332 44324
rect 45052 43148 45108 43204
rect 45388 42924 45444 42980
rect 45500 43148 45556 43204
rect 45276 42700 45332 42756
rect 46060 50540 46116 50596
rect 45948 50428 46004 50484
rect 46284 50540 46340 50596
rect 46732 50482 46788 50484
rect 46732 50430 46734 50482
rect 46734 50430 46786 50482
rect 46786 50430 46788 50482
rect 46732 50428 46788 50430
rect 46172 49026 46228 49028
rect 46172 48974 46174 49026
rect 46174 48974 46226 49026
rect 46226 48974 46228 49026
rect 46172 48972 46228 48974
rect 45836 48914 45892 48916
rect 45836 48862 45838 48914
rect 45838 48862 45890 48914
rect 45890 48862 45892 48914
rect 45836 48860 45892 48862
rect 46060 48242 46116 48244
rect 46060 48190 46062 48242
rect 46062 48190 46114 48242
rect 46114 48190 46116 48242
rect 46060 48188 46116 48190
rect 46172 47628 46228 47684
rect 46284 48076 46340 48132
rect 45948 47458 46004 47460
rect 45948 47406 45950 47458
rect 45950 47406 46002 47458
rect 46002 47406 46004 47458
rect 45948 47404 46004 47406
rect 46060 46956 46116 47012
rect 45836 46898 45892 46900
rect 45836 46846 45838 46898
rect 45838 46846 45890 46898
rect 45890 46846 45892 46898
rect 45836 46844 45892 46846
rect 45724 45218 45780 45220
rect 45724 45166 45726 45218
rect 45726 45166 45778 45218
rect 45778 45166 45780 45218
rect 45724 45164 45780 45166
rect 45836 44322 45892 44324
rect 45836 44270 45838 44322
rect 45838 44270 45890 44322
rect 45890 44270 45892 44322
rect 45836 44268 45892 44270
rect 46060 43708 46116 43764
rect 46172 43426 46228 43428
rect 46172 43374 46174 43426
rect 46174 43374 46226 43426
rect 46226 43374 46228 43426
rect 46172 43372 46228 43374
rect 45836 42978 45892 42980
rect 45836 42926 45838 42978
rect 45838 42926 45890 42978
rect 45890 42926 45892 42978
rect 45836 42924 45892 42926
rect 45724 41970 45780 41972
rect 45724 41918 45726 41970
rect 45726 41918 45778 41970
rect 45778 41918 45780 41970
rect 45724 41916 45780 41918
rect 46956 50428 47012 50484
rect 47516 51212 47572 51268
rect 47516 50652 47572 50708
rect 48188 52274 48244 52276
rect 48188 52222 48190 52274
rect 48190 52222 48242 52274
rect 48242 52222 48244 52274
rect 48188 52220 48244 52222
rect 49084 52220 49140 52276
rect 48860 52108 48916 52164
rect 48636 51436 48692 51492
rect 47292 50594 47348 50596
rect 47292 50542 47294 50594
rect 47294 50542 47346 50594
rect 47346 50542 47348 50594
rect 47292 50540 47348 50542
rect 48076 50652 48132 50708
rect 49084 50594 49140 50596
rect 49084 50542 49086 50594
rect 49086 50542 49138 50594
rect 49138 50542 49140 50594
rect 49084 50540 49140 50542
rect 46844 49810 46900 49812
rect 46844 49758 46846 49810
rect 46846 49758 46898 49810
rect 46898 49758 46900 49810
rect 46844 49756 46900 49758
rect 47180 49026 47236 49028
rect 47180 48974 47182 49026
rect 47182 48974 47234 49026
rect 47234 48974 47236 49026
rect 47180 48972 47236 48974
rect 46732 48130 46788 48132
rect 46732 48078 46734 48130
rect 46734 48078 46786 48130
rect 46786 48078 46788 48130
rect 46732 48076 46788 48078
rect 46844 47964 46900 48020
rect 47180 47458 47236 47460
rect 47180 47406 47182 47458
rect 47182 47406 47234 47458
rect 47234 47406 47236 47458
rect 47180 47404 47236 47406
rect 46956 47068 47012 47124
rect 47404 47964 47460 48020
rect 47404 47682 47460 47684
rect 47404 47630 47406 47682
rect 47406 47630 47458 47682
rect 47458 47630 47460 47682
rect 47404 47628 47460 47630
rect 46844 45164 46900 45220
rect 46620 44828 46676 44884
rect 46732 44940 46788 44996
rect 47068 45106 47124 45108
rect 47068 45054 47070 45106
rect 47070 45054 47122 45106
rect 47122 45054 47124 45106
rect 47068 45052 47124 45054
rect 47404 45052 47460 45108
rect 47180 44828 47236 44884
rect 47292 44492 47348 44548
rect 47516 44546 47572 44548
rect 47516 44494 47518 44546
rect 47518 44494 47570 44546
rect 47570 44494 47572 44546
rect 47516 44492 47572 44494
rect 46732 43762 46788 43764
rect 46732 43710 46734 43762
rect 46734 43710 46786 43762
rect 46786 43710 46788 43762
rect 46732 43708 46788 43710
rect 46508 42364 46564 42420
rect 46172 41746 46228 41748
rect 46172 41694 46174 41746
rect 46174 41694 46226 41746
rect 46226 41694 46228 41746
rect 46172 41692 46228 41694
rect 45612 40572 45668 40628
rect 46284 40908 46340 40964
rect 43372 35868 43428 35924
rect 43036 35084 43092 35140
rect 41356 34972 41412 35028
rect 42476 33346 42532 33348
rect 42476 33294 42478 33346
rect 42478 33294 42530 33346
rect 42530 33294 42532 33346
rect 42476 33292 42532 33294
rect 44044 37436 44100 37492
rect 43260 34300 43316 34356
rect 43148 33234 43204 33236
rect 43148 33182 43150 33234
rect 43150 33182 43202 33234
rect 43202 33182 43204 33234
rect 43148 33180 43204 33182
rect 43596 34690 43652 34692
rect 43596 34638 43598 34690
rect 43598 34638 43650 34690
rect 43650 34638 43652 34690
rect 43596 34636 43652 34638
rect 43932 34636 43988 34692
rect 43932 33628 43988 33684
rect 43148 32956 43204 33012
rect 42700 32172 42756 32228
rect 41692 31218 41748 31220
rect 41692 31166 41694 31218
rect 41694 31166 41746 31218
rect 41746 31166 41748 31218
rect 41692 31164 41748 31166
rect 41916 31218 41972 31220
rect 41916 31166 41918 31218
rect 41918 31166 41970 31218
rect 41970 31166 41972 31218
rect 41916 31164 41972 31166
rect 39788 30940 39844 30996
rect 41356 30994 41412 30996
rect 41356 30942 41358 30994
rect 41358 30942 41410 30994
rect 41410 30942 41412 30994
rect 41356 30940 41412 30942
rect 40348 30828 40404 30884
rect 39676 30380 39732 30436
rect 37324 29596 37380 29652
rect 41020 30882 41076 30884
rect 41020 30830 41022 30882
rect 41022 30830 41074 30882
rect 41074 30830 41076 30882
rect 41020 30828 41076 30830
rect 38444 29650 38500 29652
rect 38444 29598 38446 29650
rect 38446 29598 38498 29650
rect 38498 29598 38500 29650
rect 38444 29596 38500 29598
rect 38556 29932 38612 29988
rect 33740 29426 33796 29428
rect 33740 29374 33742 29426
rect 33742 29374 33794 29426
rect 33794 29374 33796 29426
rect 33740 29372 33796 29374
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 33964 28754 34020 28756
rect 33964 28702 33966 28754
rect 33966 28702 34018 28754
rect 34018 28702 34020 28754
rect 33964 28700 34020 28702
rect 34972 28588 35028 28644
rect 32956 28418 33012 28420
rect 32956 28366 32958 28418
rect 32958 28366 33010 28418
rect 33010 28366 33012 28418
rect 32956 28364 33012 28366
rect 33964 28028 34020 28084
rect 31724 27132 31780 27188
rect 32284 27132 32340 27188
rect 29372 26236 29428 26292
rect 29148 25564 29204 25620
rect 28588 25506 28644 25508
rect 28588 25454 28590 25506
rect 28590 25454 28642 25506
rect 28642 25454 28644 25506
rect 28588 25452 28644 25454
rect 28252 25116 28308 25172
rect 28364 25340 28420 25396
rect 28476 25116 28532 25172
rect 28700 24834 28756 24836
rect 28700 24782 28702 24834
rect 28702 24782 28754 24834
rect 28754 24782 28756 24834
rect 28700 24780 28756 24782
rect 28364 23212 28420 23268
rect 28140 23100 28196 23156
rect 27692 20636 27748 20692
rect 27580 20300 27636 20356
rect 27468 20130 27524 20132
rect 27468 20078 27470 20130
rect 27470 20078 27522 20130
rect 27522 20078 27524 20130
rect 27468 20076 27524 20078
rect 27580 19852 27636 19908
rect 27468 18844 27524 18900
rect 27692 18508 27748 18564
rect 27692 18338 27748 18340
rect 27692 18286 27694 18338
rect 27694 18286 27746 18338
rect 27746 18286 27748 18338
rect 27692 18284 27748 18286
rect 27692 17276 27748 17332
rect 27468 16716 27524 16772
rect 27356 12460 27412 12516
rect 27356 12012 27412 12068
rect 27580 16156 27636 16212
rect 27804 17164 27860 17220
rect 28140 20130 28196 20132
rect 28140 20078 28142 20130
rect 28142 20078 28194 20130
rect 28194 20078 28196 20130
rect 28140 20076 28196 20078
rect 28476 20802 28532 20804
rect 28476 20750 28478 20802
rect 28478 20750 28530 20802
rect 28530 20750 28532 20802
rect 28476 20748 28532 20750
rect 28364 20300 28420 20356
rect 29260 25394 29316 25396
rect 29260 25342 29262 25394
rect 29262 25342 29314 25394
rect 29314 25342 29316 25394
rect 29260 25340 29316 25342
rect 30380 26290 30436 26292
rect 30380 26238 30382 26290
rect 30382 26238 30434 26290
rect 30434 26238 30436 26290
rect 30380 26236 30436 26238
rect 30268 25900 30324 25956
rect 29708 25788 29764 25844
rect 29596 25116 29652 25172
rect 28588 20130 28644 20132
rect 28588 20078 28590 20130
rect 28590 20078 28642 20130
rect 28642 20078 28644 20130
rect 28588 20076 28644 20078
rect 28140 19516 28196 19572
rect 28476 19180 28532 19236
rect 28588 18732 28644 18788
rect 28252 17890 28308 17892
rect 28252 17838 28254 17890
rect 28254 17838 28306 17890
rect 28306 17838 28308 17890
rect 28252 17836 28308 17838
rect 28028 16940 28084 16996
rect 28364 17164 28420 17220
rect 27916 16156 27972 16212
rect 27804 16098 27860 16100
rect 27804 16046 27806 16098
rect 27806 16046 27858 16098
rect 27858 16046 27860 16098
rect 27804 16044 27860 16046
rect 27580 15372 27636 15428
rect 27692 15596 27748 15652
rect 27916 15260 27972 15316
rect 27804 14418 27860 14420
rect 27804 14366 27806 14418
rect 27806 14366 27858 14418
rect 27858 14366 27860 14418
rect 27804 14364 27860 14366
rect 27692 13356 27748 13412
rect 27244 11676 27300 11732
rect 27692 12908 27748 12964
rect 27804 13692 27860 13748
rect 28140 15538 28196 15540
rect 28140 15486 28142 15538
rect 28142 15486 28194 15538
rect 28194 15486 28196 15538
rect 28140 15484 28196 15486
rect 28924 19852 28980 19908
rect 28812 18396 28868 18452
rect 28700 16492 28756 16548
rect 29484 23266 29540 23268
rect 29484 23214 29486 23266
rect 29486 23214 29538 23266
rect 29538 23214 29540 23266
rect 29484 23212 29540 23214
rect 29260 22258 29316 22260
rect 29260 22206 29262 22258
rect 29262 22206 29314 22258
rect 29314 22206 29316 22258
rect 29260 22204 29316 22206
rect 29148 21420 29204 21476
rect 29148 20860 29204 20916
rect 29932 25564 29988 25620
rect 30044 25506 30100 25508
rect 30044 25454 30046 25506
rect 30046 25454 30098 25506
rect 30098 25454 30100 25506
rect 30044 25452 30100 25454
rect 30156 24780 30212 24836
rect 29932 22540 29988 22596
rect 29820 21644 29876 21700
rect 29820 20748 29876 20804
rect 29148 19516 29204 19572
rect 29260 18732 29316 18788
rect 29484 18620 29540 18676
rect 30044 19964 30100 20020
rect 29932 19516 29988 19572
rect 29708 17724 29764 17780
rect 28588 15596 28644 15652
rect 28140 14924 28196 14980
rect 27580 12236 27636 12292
rect 27244 11452 27300 11508
rect 26908 10498 26964 10500
rect 26908 10446 26910 10498
rect 26910 10446 26962 10498
rect 26962 10446 26964 10498
rect 26908 10444 26964 10446
rect 27692 12684 27748 12740
rect 27916 13020 27972 13076
rect 27804 12124 27860 12180
rect 27580 11170 27636 11172
rect 27580 11118 27582 11170
rect 27582 11118 27634 11170
rect 27634 11118 27636 11170
rect 27580 11116 27636 11118
rect 26796 9266 26852 9268
rect 26796 9214 26798 9266
rect 26798 9214 26850 9266
rect 26850 9214 26852 9266
rect 26796 9212 26852 9214
rect 26684 8764 26740 8820
rect 26796 8652 26852 8708
rect 26572 6860 26628 6916
rect 27580 9996 27636 10052
rect 27468 9884 27524 9940
rect 27356 9324 27412 9380
rect 28140 14252 28196 14308
rect 28140 12962 28196 12964
rect 28140 12910 28142 12962
rect 28142 12910 28194 12962
rect 28194 12910 28196 12962
rect 28140 12908 28196 12910
rect 28140 12572 28196 12628
rect 28364 15148 28420 15204
rect 28924 15932 28980 15988
rect 29036 15820 29092 15876
rect 28588 13634 28644 13636
rect 28588 13582 28590 13634
rect 28590 13582 28642 13634
rect 28642 13582 28644 13634
rect 28588 13580 28644 13582
rect 28476 13132 28532 13188
rect 28924 13356 28980 13412
rect 28700 11900 28756 11956
rect 28812 11788 28868 11844
rect 28476 11676 28532 11732
rect 28700 11452 28756 11508
rect 27692 9826 27748 9828
rect 27692 9774 27694 9826
rect 27694 9774 27746 9826
rect 27746 9774 27748 9826
rect 27692 9772 27748 9774
rect 28364 9772 28420 9828
rect 27916 9266 27972 9268
rect 27916 9214 27918 9266
rect 27918 9214 27970 9266
rect 27970 9214 27972 9266
rect 27916 9212 27972 9214
rect 28812 11340 28868 11396
rect 29260 16492 29316 16548
rect 29708 16716 29764 16772
rect 29708 16210 29764 16212
rect 29708 16158 29710 16210
rect 29710 16158 29762 16210
rect 29762 16158 29764 16210
rect 29708 16156 29764 16158
rect 29484 15932 29540 15988
rect 29372 15484 29428 15540
rect 29596 15314 29652 15316
rect 29596 15262 29598 15314
rect 29598 15262 29650 15314
rect 29650 15262 29652 15314
rect 29596 15260 29652 15262
rect 29820 15820 29876 15876
rect 29372 14364 29428 14420
rect 29148 13580 29204 13636
rect 29372 13692 29428 13748
rect 29484 13804 29540 13860
rect 29932 13580 29988 13636
rect 29596 13468 29652 13524
rect 30380 19516 30436 19572
rect 30716 26012 30772 26068
rect 31052 26012 31108 26068
rect 31276 25900 31332 25956
rect 32060 25676 32116 25732
rect 31836 25228 31892 25284
rect 30604 25116 30660 25172
rect 30604 24946 30660 24948
rect 30604 24894 30606 24946
rect 30606 24894 30658 24946
rect 30658 24894 30660 24946
rect 30604 24892 30660 24894
rect 31164 24780 31220 24836
rect 31164 24050 31220 24052
rect 31164 23998 31166 24050
rect 31166 23998 31218 24050
rect 31218 23998 31220 24050
rect 31164 23996 31220 23998
rect 31836 24722 31892 24724
rect 31836 24670 31838 24722
rect 31838 24670 31890 24722
rect 31890 24670 31892 24722
rect 31836 24668 31892 24670
rect 31388 23548 31444 23604
rect 31948 23660 32004 23716
rect 31276 23154 31332 23156
rect 31276 23102 31278 23154
rect 31278 23102 31330 23154
rect 31330 23102 31332 23154
rect 31276 23100 31332 23102
rect 30604 21474 30660 21476
rect 30604 21422 30606 21474
rect 30606 21422 30658 21474
rect 30658 21422 30660 21474
rect 30604 21420 30660 21422
rect 30492 18562 30548 18564
rect 30492 18510 30494 18562
rect 30494 18510 30546 18562
rect 30546 18510 30548 18562
rect 30492 18508 30548 18510
rect 30716 20242 30772 20244
rect 30716 20190 30718 20242
rect 30718 20190 30770 20242
rect 30770 20190 30772 20242
rect 30716 20188 30772 20190
rect 31164 21756 31220 21812
rect 31052 21698 31108 21700
rect 31052 21646 31054 21698
rect 31054 21646 31106 21698
rect 31106 21646 31108 21698
rect 31052 21644 31108 21646
rect 31500 22482 31556 22484
rect 31500 22430 31502 22482
rect 31502 22430 31554 22482
rect 31554 22430 31556 22482
rect 31500 22428 31556 22430
rect 32172 25618 32228 25620
rect 32172 25566 32174 25618
rect 32174 25566 32226 25618
rect 32226 25566 32228 25618
rect 32172 25564 32228 25566
rect 32060 23100 32116 23156
rect 35644 28588 35700 28644
rect 35532 28476 35588 28532
rect 35532 27634 35588 27636
rect 35532 27582 35534 27634
rect 35534 27582 35586 27634
rect 35586 27582 35588 27634
rect 35532 27580 35588 27582
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35756 27468 35812 27524
rect 35756 27186 35812 27188
rect 35756 27134 35758 27186
rect 35758 27134 35810 27186
rect 35810 27134 35812 27186
rect 35756 27132 35812 27134
rect 37324 28700 37380 28756
rect 37212 28642 37268 28644
rect 37212 28590 37214 28642
rect 37214 28590 37266 28642
rect 37266 28590 37268 28642
rect 37212 28588 37268 28590
rect 37100 28530 37156 28532
rect 37100 28478 37102 28530
rect 37102 28478 37154 28530
rect 37154 28478 37156 28530
rect 37100 28476 37156 28478
rect 36876 27916 36932 27972
rect 36428 27132 36484 27188
rect 37100 27186 37156 27188
rect 37100 27134 37102 27186
rect 37102 27134 37154 27186
rect 37154 27134 37156 27186
rect 37100 27132 37156 27134
rect 34972 27020 35028 27076
rect 36988 27074 37044 27076
rect 36988 27022 36990 27074
rect 36990 27022 37042 27074
rect 37042 27022 37044 27074
rect 36988 27020 37044 27022
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35196 25564 35252 25620
rect 36092 25618 36148 25620
rect 36092 25566 36094 25618
rect 36094 25566 36146 25618
rect 36146 25566 36148 25618
rect 36092 25564 36148 25566
rect 33180 24722 33236 24724
rect 33180 24670 33182 24722
rect 33182 24670 33234 24722
rect 33234 24670 33236 24722
rect 33180 24668 33236 24670
rect 33404 23938 33460 23940
rect 33404 23886 33406 23938
rect 33406 23886 33458 23938
rect 33458 23886 33460 23938
rect 33404 23884 33460 23886
rect 33852 24668 33908 24724
rect 33740 23884 33796 23940
rect 32508 23154 32564 23156
rect 32508 23102 32510 23154
rect 32510 23102 32562 23154
rect 32562 23102 32564 23154
rect 32508 23100 32564 23102
rect 33628 23154 33684 23156
rect 33628 23102 33630 23154
rect 33630 23102 33682 23154
rect 33682 23102 33684 23154
rect 33628 23100 33684 23102
rect 33516 22988 33572 23044
rect 32396 22428 32452 22484
rect 31388 21756 31444 21812
rect 32172 21756 32228 21812
rect 31164 21196 31220 21252
rect 30940 20748 30996 20804
rect 31052 20636 31108 20692
rect 31612 21196 31668 21252
rect 32508 21362 32564 21364
rect 32508 21310 32510 21362
rect 32510 21310 32562 21362
rect 32562 21310 32564 21362
rect 32508 21308 32564 21310
rect 32396 20972 32452 21028
rect 31948 20748 32004 20804
rect 31724 20242 31780 20244
rect 31724 20190 31726 20242
rect 31726 20190 31778 20242
rect 31778 20190 31780 20242
rect 31724 20188 31780 20190
rect 32284 20748 32340 20804
rect 32172 20412 32228 20468
rect 30604 18172 30660 18228
rect 30380 16156 30436 16212
rect 30492 16940 30548 16996
rect 30492 15036 30548 15092
rect 30492 14252 30548 14308
rect 30492 14028 30548 14084
rect 31276 19292 31332 19348
rect 30940 19180 30996 19236
rect 31948 19628 32004 19684
rect 31612 19292 31668 19348
rect 31052 16940 31108 16996
rect 31612 19010 31668 19012
rect 31612 18958 31614 19010
rect 31614 18958 31666 19010
rect 31666 18958 31668 19010
rect 31612 18956 31668 18958
rect 32732 19346 32788 19348
rect 32732 19294 32734 19346
rect 32734 19294 32786 19346
rect 32786 19294 32788 19346
rect 32732 19292 32788 19294
rect 32620 17778 32676 17780
rect 32620 17726 32622 17778
rect 32622 17726 32674 17778
rect 32674 17726 32676 17778
rect 32620 17724 32676 17726
rect 31164 16828 31220 16884
rect 30828 15874 30884 15876
rect 30828 15822 30830 15874
rect 30830 15822 30882 15874
rect 30882 15822 30884 15874
rect 30828 15820 30884 15822
rect 31276 15260 31332 15316
rect 29260 12066 29316 12068
rect 29260 12014 29262 12066
rect 29262 12014 29314 12066
rect 29314 12014 29316 12066
rect 29260 12012 29316 12014
rect 29596 11452 29652 11508
rect 30492 13858 30548 13860
rect 30492 13806 30494 13858
rect 30494 13806 30546 13858
rect 30546 13806 30548 13858
rect 30492 13804 30548 13806
rect 30604 13746 30660 13748
rect 30604 13694 30606 13746
rect 30606 13694 30658 13746
rect 30658 13694 30660 13746
rect 30604 13692 30660 13694
rect 30044 12236 30100 12292
rect 30268 12290 30324 12292
rect 30268 12238 30270 12290
rect 30270 12238 30322 12290
rect 30322 12238 30324 12290
rect 30268 12236 30324 12238
rect 29932 12178 29988 12180
rect 29932 12126 29934 12178
rect 29934 12126 29986 12178
rect 29986 12126 29988 12178
rect 29932 12124 29988 12126
rect 30492 12178 30548 12180
rect 30492 12126 30494 12178
rect 30494 12126 30546 12178
rect 30546 12126 30548 12178
rect 30492 12124 30548 12126
rect 29708 12012 29764 12068
rect 29260 11228 29316 11284
rect 29148 10444 29204 10500
rect 27804 8876 27860 8932
rect 26460 6636 26516 6692
rect 26236 6524 26292 6580
rect 26348 6300 26404 6356
rect 25900 5906 25956 5908
rect 25900 5854 25902 5906
rect 25902 5854 25954 5906
rect 25954 5854 25956 5906
rect 25900 5852 25956 5854
rect 26236 6188 26292 6244
rect 25788 5292 25844 5348
rect 25564 4396 25620 4452
rect 26796 6412 26852 6468
rect 26684 5964 26740 6020
rect 27244 8034 27300 8036
rect 27244 7982 27246 8034
rect 27246 7982 27298 8034
rect 27298 7982 27300 8034
rect 27244 7980 27300 7982
rect 27580 8146 27636 8148
rect 27580 8094 27582 8146
rect 27582 8094 27634 8146
rect 27634 8094 27636 8146
rect 27580 8092 27636 8094
rect 28364 8146 28420 8148
rect 28364 8094 28366 8146
rect 28366 8094 28418 8146
rect 28418 8094 28420 8146
rect 28364 8092 28420 8094
rect 28476 7980 28532 8036
rect 29148 9826 29204 9828
rect 29148 9774 29150 9826
rect 29150 9774 29202 9826
rect 29202 9774 29204 9826
rect 29148 9772 29204 9774
rect 31052 13858 31108 13860
rect 31052 13806 31054 13858
rect 31054 13806 31106 13858
rect 31106 13806 31108 13858
rect 31052 13804 31108 13806
rect 31276 14028 31332 14084
rect 31724 17554 31780 17556
rect 31724 17502 31726 17554
rect 31726 17502 31778 17554
rect 31778 17502 31780 17554
rect 31724 17500 31780 17502
rect 31836 16604 31892 16660
rect 31612 15596 31668 15652
rect 31724 15820 31780 15876
rect 31500 14812 31556 14868
rect 31052 12738 31108 12740
rect 31052 12686 31054 12738
rect 31054 12686 31106 12738
rect 31106 12686 31108 12738
rect 31052 12684 31108 12686
rect 31052 12460 31108 12516
rect 30940 12348 30996 12404
rect 31836 14812 31892 14868
rect 31388 12684 31444 12740
rect 31500 12572 31556 12628
rect 31388 12348 31444 12404
rect 31052 12124 31108 12180
rect 31164 11954 31220 11956
rect 31164 11902 31166 11954
rect 31166 11902 31218 11954
rect 31218 11902 31220 11954
rect 31164 11900 31220 11902
rect 30156 11676 30212 11732
rect 29932 11228 29988 11284
rect 30156 10834 30212 10836
rect 30156 10782 30158 10834
rect 30158 10782 30210 10834
rect 30210 10782 30212 10834
rect 30156 10780 30212 10782
rect 30044 10498 30100 10500
rect 30044 10446 30046 10498
rect 30046 10446 30098 10498
rect 30098 10446 30100 10498
rect 30044 10444 30100 10446
rect 29932 10332 29988 10388
rect 30268 9996 30324 10052
rect 29596 9436 29652 9492
rect 29372 9212 29428 9268
rect 29260 9154 29316 9156
rect 29260 9102 29262 9154
rect 29262 9102 29314 9154
rect 29314 9102 29316 9154
rect 29260 9100 29316 9102
rect 29708 9154 29764 9156
rect 29708 9102 29710 9154
rect 29710 9102 29762 9154
rect 29762 9102 29764 9154
rect 29708 9100 29764 9102
rect 28252 7698 28308 7700
rect 28252 7646 28254 7698
rect 28254 7646 28306 7698
rect 28306 7646 28308 7698
rect 28252 7644 28308 7646
rect 29596 8034 29652 8036
rect 29596 7982 29598 8034
rect 29598 7982 29650 8034
rect 29650 7982 29652 8034
rect 29596 7980 29652 7982
rect 29036 7644 29092 7700
rect 27580 7420 27636 7476
rect 28028 7308 28084 7364
rect 26908 5964 26964 6020
rect 27244 6972 27300 7028
rect 27468 6076 27524 6132
rect 27692 5964 27748 6020
rect 26908 5516 26964 5572
rect 27020 5180 27076 5236
rect 25004 2828 25060 2884
rect 16604 2604 16660 2660
rect 28140 6578 28196 6580
rect 28140 6526 28142 6578
rect 28142 6526 28194 6578
rect 28194 6526 28196 6578
rect 28140 6524 28196 6526
rect 28812 6748 28868 6804
rect 28476 6690 28532 6692
rect 28476 6638 28478 6690
rect 28478 6638 28530 6690
rect 28530 6638 28532 6690
rect 28476 6636 28532 6638
rect 28364 6524 28420 6580
rect 28812 6412 28868 6468
rect 28140 5906 28196 5908
rect 28140 5854 28142 5906
rect 28142 5854 28194 5906
rect 28194 5854 28196 5906
rect 28140 5852 28196 5854
rect 29708 7420 29764 7476
rect 29260 6802 29316 6804
rect 29260 6750 29262 6802
rect 29262 6750 29314 6802
rect 29314 6750 29316 6802
rect 29260 6748 29316 6750
rect 29036 5964 29092 6020
rect 29820 6748 29876 6804
rect 30268 8428 30324 8484
rect 30044 8146 30100 8148
rect 30044 8094 30046 8146
rect 30046 8094 30098 8146
rect 30098 8094 30100 8146
rect 30044 8092 30100 8094
rect 30380 8146 30436 8148
rect 30380 8094 30382 8146
rect 30382 8094 30434 8146
rect 30434 8094 30436 8146
rect 30380 8092 30436 8094
rect 30156 8034 30212 8036
rect 30156 7982 30158 8034
rect 30158 7982 30210 8034
rect 30210 7982 30212 8034
rect 30156 7980 30212 7982
rect 29932 6130 29988 6132
rect 29932 6078 29934 6130
rect 29934 6078 29986 6130
rect 29986 6078 29988 6130
rect 29932 6076 29988 6078
rect 29372 5852 29428 5908
rect 27804 5292 27860 5348
rect 28476 5404 28532 5460
rect 28476 5122 28532 5124
rect 28476 5070 28478 5122
rect 28478 5070 28530 5122
rect 28530 5070 28532 5122
rect 28476 5068 28532 5070
rect 28812 5292 28868 5348
rect 28140 4956 28196 5012
rect 28140 4732 28196 4788
rect 29148 5180 29204 5236
rect 30380 5234 30436 5236
rect 30380 5182 30382 5234
rect 30382 5182 30434 5234
rect 30434 5182 30436 5234
rect 30380 5180 30436 5182
rect 29484 5068 29540 5124
rect 29708 5010 29764 5012
rect 29708 4958 29710 5010
rect 29710 4958 29762 5010
rect 29762 4958 29764 5010
rect 29708 4956 29764 4958
rect 30380 4562 30436 4564
rect 30380 4510 30382 4562
rect 30382 4510 30434 4562
rect 30434 4510 30436 4562
rect 30380 4508 30436 4510
rect 28812 3666 28868 3668
rect 28812 3614 28814 3666
rect 28814 3614 28866 3666
rect 28866 3614 28868 3666
rect 28812 3612 28868 3614
rect 27132 2604 27188 2660
rect 28924 3388 28980 3444
rect 30044 3388 30100 3444
rect 31388 11506 31444 11508
rect 31388 11454 31390 11506
rect 31390 11454 31442 11506
rect 31442 11454 31444 11506
rect 31388 11452 31444 11454
rect 31052 11394 31108 11396
rect 31052 11342 31054 11394
rect 31054 11342 31106 11394
rect 31106 11342 31108 11394
rect 31052 11340 31108 11342
rect 30940 11282 30996 11284
rect 30940 11230 30942 11282
rect 30942 11230 30994 11282
rect 30994 11230 30996 11282
rect 30940 11228 30996 11230
rect 30604 10668 30660 10724
rect 31276 10498 31332 10500
rect 31276 10446 31278 10498
rect 31278 10446 31330 10498
rect 31330 10446 31332 10498
rect 31276 10444 31332 10446
rect 30604 6130 30660 6132
rect 30604 6078 30606 6130
rect 30606 6078 30658 6130
rect 30658 6078 30660 6130
rect 30604 6076 30660 6078
rect 30716 4620 30772 4676
rect 33292 20188 33348 20244
rect 33068 19292 33124 19348
rect 33516 22428 33572 22484
rect 33964 24556 34020 24612
rect 33852 21868 33908 21924
rect 33516 21196 33572 21252
rect 33516 20412 33572 20468
rect 33628 20130 33684 20132
rect 33628 20078 33630 20130
rect 33630 20078 33682 20130
rect 33682 20078 33684 20130
rect 33628 20076 33684 20078
rect 33628 19740 33684 19796
rect 33852 21532 33908 21588
rect 33852 20524 33908 20580
rect 34972 24556 35028 24612
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 34860 23100 34916 23156
rect 34300 23042 34356 23044
rect 34300 22990 34302 23042
rect 34302 22990 34354 23042
rect 34354 22990 34356 23042
rect 34300 22988 34356 22990
rect 36204 25282 36260 25284
rect 36204 25230 36206 25282
rect 36206 25230 36258 25282
rect 36258 25230 36260 25282
rect 36204 25228 36260 25230
rect 36988 25282 37044 25284
rect 36988 25230 36990 25282
rect 36990 25230 37042 25282
rect 37042 25230 37044 25282
rect 36988 25228 37044 25230
rect 35756 23660 35812 23716
rect 35196 23100 35252 23156
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 34524 22316 34580 22372
rect 33740 19628 33796 19684
rect 33404 17948 33460 18004
rect 33404 17554 33460 17556
rect 33404 17502 33406 17554
rect 33406 17502 33458 17554
rect 33458 17502 33460 17554
rect 33404 17500 33460 17502
rect 34972 21756 35028 21812
rect 36876 24556 36932 24612
rect 36092 23884 36148 23940
rect 35980 23100 36036 23156
rect 36988 23660 37044 23716
rect 36204 22482 36260 22484
rect 36204 22430 36206 22482
rect 36206 22430 36258 22482
rect 36258 22430 36260 22482
rect 36204 22428 36260 22430
rect 35980 22370 36036 22372
rect 35980 22318 35982 22370
rect 35982 22318 36034 22370
rect 36034 22318 36036 22370
rect 35980 22316 36036 22318
rect 36204 22204 36260 22260
rect 34636 21474 34692 21476
rect 34636 21422 34638 21474
rect 34638 21422 34690 21474
rect 34690 21422 34692 21474
rect 34636 21420 34692 21422
rect 35084 21532 35140 21588
rect 35644 21532 35700 21588
rect 35084 21308 35140 21364
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 34748 20860 34804 20916
rect 34076 20076 34132 20132
rect 34524 19964 34580 20020
rect 34300 19906 34356 19908
rect 34300 19854 34302 19906
rect 34302 19854 34354 19906
rect 34354 19854 34356 19906
rect 34300 19852 34356 19854
rect 33964 19010 34020 19012
rect 33964 18958 33966 19010
rect 33966 18958 34018 19010
rect 34018 18958 34020 19010
rect 33964 18956 34020 18958
rect 34524 18956 34580 19012
rect 34748 20300 34804 20356
rect 35868 20914 35924 20916
rect 35868 20862 35870 20914
rect 35870 20862 35922 20914
rect 35922 20862 35924 20914
rect 35868 20860 35924 20862
rect 36316 21532 36372 21588
rect 34972 20076 35028 20132
rect 35980 19740 36036 19796
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 34300 17948 34356 18004
rect 34300 17666 34356 17668
rect 34300 17614 34302 17666
rect 34302 17614 34354 17666
rect 34354 17614 34356 17666
rect 34300 17612 34356 17614
rect 34076 17500 34132 17556
rect 33404 16156 33460 16212
rect 32956 15932 33012 15988
rect 32956 15314 33012 15316
rect 32956 15262 32958 15314
rect 32958 15262 33010 15314
rect 33010 15262 33012 15314
rect 32956 15260 33012 15262
rect 32172 14476 32228 14532
rect 32396 14588 32452 14644
rect 31948 14364 32004 14420
rect 32284 13692 32340 13748
rect 31836 10722 31892 10724
rect 31836 10670 31838 10722
rect 31838 10670 31890 10722
rect 31890 10670 31892 10722
rect 31836 10668 31892 10670
rect 31724 9996 31780 10052
rect 31500 9212 31556 9268
rect 31612 9548 31668 9604
rect 31724 8204 31780 8260
rect 32060 8258 32116 8260
rect 32060 8206 32062 8258
rect 32062 8206 32114 8258
rect 32114 8206 32116 8258
rect 32060 8204 32116 8206
rect 33516 16098 33572 16100
rect 33516 16046 33518 16098
rect 33518 16046 33570 16098
rect 33570 16046 33572 16098
rect 33516 16044 33572 16046
rect 33628 15986 33684 15988
rect 33628 15934 33630 15986
rect 33630 15934 33682 15986
rect 33682 15934 33684 15986
rect 33628 15932 33684 15934
rect 33180 15874 33236 15876
rect 33180 15822 33182 15874
rect 33182 15822 33234 15874
rect 33234 15822 33236 15874
rect 33180 15820 33236 15822
rect 33404 15148 33460 15204
rect 33404 14924 33460 14980
rect 33292 14140 33348 14196
rect 32508 13580 32564 13636
rect 33516 14700 33572 14756
rect 33964 16156 34020 16212
rect 34748 17836 34804 17892
rect 34524 17500 34580 17556
rect 34412 16882 34468 16884
rect 34412 16830 34414 16882
rect 34414 16830 34466 16882
rect 34466 16830 34468 16882
rect 34412 16828 34468 16830
rect 34412 16156 34468 16212
rect 34300 16098 34356 16100
rect 34300 16046 34302 16098
rect 34302 16046 34354 16098
rect 34354 16046 34356 16098
rect 34300 16044 34356 16046
rect 34076 15932 34132 15988
rect 34076 15484 34132 15540
rect 33740 14924 33796 14980
rect 33964 15202 34020 15204
rect 33964 15150 33966 15202
rect 33966 15150 34018 15202
rect 34018 15150 34020 15202
rect 33964 15148 34020 15150
rect 33628 14588 33684 14644
rect 33628 14418 33684 14420
rect 33628 14366 33630 14418
rect 33630 14366 33682 14418
rect 33682 14366 33684 14418
rect 33628 14364 33684 14366
rect 33628 13858 33684 13860
rect 33628 13806 33630 13858
rect 33630 13806 33682 13858
rect 33682 13806 33684 13858
rect 33628 13804 33684 13806
rect 33852 13746 33908 13748
rect 33852 13694 33854 13746
rect 33854 13694 33906 13746
rect 33906 13694 33908 13746
rect 33852 13692 33908 13694
rect 32956 11564 33012 11620
rect 33740 11564 33796 11620
rect 33516 11340 33572 11396
rect 33740 10892 33796 10948
rect 33628 10668 33684 10724
rect 32956 10220 33012 10276
rect 32620 9996 32676 10052
rect 32396 9212 32452 9268
rect 32508 8930 32564 8932
rect 32508 8878 32510 8930
rect 32510 8878 32562 8930
rect 32562 8878 32564 8930
rect 32508 8876 32564 8878
rect 32060 7980 32116 8036
rect 31948 7532 32004 7588
rect 31612 6690 31668 6692
rect 31612 6638 31614 6690
rect 31614 6638 31666 6690
rect 31666 6638 31668 6690
rect 31612 6636 31668 6638
rect 32508 7586 32564 7588
rect 32508 7534 32510 7586
rect 32510 7534 32562 7586
rect 32562 7534 32564 7586
rect 32508 7532 32564 7534
rect 32732 7980 32788 8036
rect 33068 8146 33124 8148
rect 33068 8094 33070 8146
rect 33070 8094 33122 8146
rect 33122 8094 33124 8146
rect 33068 8092 33124 8094
rect 33180 8034 33236 8036
rect 33180 7982 33182 8034
rect 33182 7982 33234 8034
rect 33234 7982 33236 8034
rect 33180 7980 33236 7982
rect 33516 7532 33572 7588
rect 32620 6748 32676 6804
rect 32956 6636 33012 6692
rect 32508 6524 32564 6580
rect 32172 6300 32228 6356
rect 31612 5180 31668 5236
rect 32732 5234 32788 5236
rect 32732 5182 32734 5234
rect 32734 5182 32786 5234
rect 32786 5182 32788 5234
rect 32732 5180 32788 5182
rect 30604 4338 30660 4340
rect 30604 4286 30606 4338
rect 30606 4286 30658 4338
rect 30658 4286 30660 4338
rect 30604 4284 30660 4286
rect 32284 4844 32340 4900
rect 31836 4338 31892 4340
rect 31836 4286 31838 4338
rect 31838 4286 31890 4338
rect 31890 4286 31892 4338
rect 31836 4284 31892 4286
rect 33068 4562 33124 4564
rect 33068 4510 33070 4562
rect 33070 4510 33122 4562
rect 33122 4510 33124 4562
rect 33068 4508 33124 4510
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35420 17724 35476 17780
rect 35756 17836 35812 17892
rect 36540 20018 36596 20020
rect 36540 19966 36542 20018
rect 36542 19966 36594 20018
rect 36594 19966 36596 20018
rect 36540 19964 36596 19966
rect 36428 18844 36484 18900
rect 35980 17724 36036 17780
rect 35532 17612 35588 17668
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 36092 16940 36148 16996
rect 36428 16882 36484 16884
rect 36428 16830 36430 16882
rect 36430 16830 36482 16882
rect 36482 16830 36484 16882
rect 36428 16828 36484 16830
rect 36316 16604 36372 16660
rect 35980 16210 36036 16212
rect 35980 16158 35982 16210
rect 35982 16158 36034 16210
rect 36034 16158 36036 16210
rect 35980 16156 36036 16158
rect 35196 16044 35252 16100
rect 35756 15986 35812 15988
rect 35756 15934 35758 15986
rect 35758 15934 35810 15986
rect 35810 15934 35812 15986
rect 35756 15932 35812 15934
rect 35084 15484 35140 15540
rect 36092 15260 36148 15316
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35084 14530 35140 14532
rect 35084 14478 35086 14530
rect 35086 14478 35138 14530
rect 35138 14478 35140 14530
rect 35084 14476 35140 14478
rect 34972 14364 35028 14420
rect 35084 13858 35140 13860
rect 35084 13806 35086 13858
rect 35086 13806 35138 13858
rect 35138 13806 35140 13858
rect 35084 13804 35140 13806
rect 35532 14588 35588 14644
rect 35308 14140 35364 14196
rect 35196 13692 35252 13748
rect 34636 13634 34692 13636
rect 34636 13582 34638 13634
rect 34638 13582 34690 13634
rect 34690 13582 34692 13634
rect 34636 13580 34692 13582
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 36316 14642 36372 14644
rect 36316 14590 36318 14642
rect 36318 14590 36370 14642
rect 36370 14590 36372 14642
rect 36316 14588 36372 14590
rect 35196 12402 35252 12404
rect 35196 12350 35198 12402
rect 35198 12350 35250 12402
rect 35250 12350 35252 12402
rect 35196 12348 35252 12350
rect 35756 12348 35812 12404
rect 36428 12348 36484 12404
rect 34748 12178 34804 12180
rect 34748 12126 34750 12178
rect 34750 12126 34802 12178
rect 34802 12126 34804 12178
rect 34748 12124 34804 12126
rect 35980 12178 36036 12180
rect 35980 12126 35982 12178
rect 35982 12126 36034 12178
rect 36034 12126 36036 12178
rect 35980 12124 36036 12126
rect 35868 11900 35924 11956
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 34076 11394 34132 11396
rect 34076 11342 34078 11394
rect 34078 11342 34130 11394
rect 34130 11342 34132 11394
rect 34076 11340 34132 11342
rect 34188 11564 34244 11620
rect 34076 10332 34132 10388
rect 34300 11452 34356 11508
rect 34748 11452 34804 11508
rect 34636 11340 34692 11396
rect 34524 11282 34580 11284
rect 34524 11230 34526 11282
rect 34526 11230 34578 11282
rect 34578 11230 34580 11282
rect 34524 11228 34580 11230
rect 35196 11452 35252 11508
rect 35308 11394 35364 11396
rect 35308 11342 35310 11394
rect 35310 11342 35362 11394
rect 35362 11342 35364 11394
rect 35308 11340 35364 11342
rect 34972 10722 35028 10724
rect 34972 10670 34974 10722
rect 34974 10670 35026 10722
rect 35026 10670 35028 10722
rect 34972 10668 35028 10670
rect 34412 7586 34468 7588
rect 34412 7534 34414 7586
rect 34414 7534 34466 7586
rect 34466 7534 34468 7586
rect 34412 7532 34468 7534
rect 33964 6690 34020 6692
rect 33964 6638 33966 6690
rect 33966 6638 34018 6690
rect 34018 6638 34020 6690
rect 33964 6636 34020 6638
rect 35420 10332 35476 10388
rect 36092 11676 36148 11732
rect 37548 28588 37604 28644
rect 37436 27580 37492 27636
rect 38220 28642 38276 28644
rect 38220 28590 38222 28642
rect 38222 28590 38274 28642
rect 38274 28590 38276 28642
rect 38220 28588 38276 28590
rect 38332 28476 38388 28532
rect 39228 29986 39284 29988
rect 39228 29934 39230 29986
rect 39230 29934 39282 29986
rect 39282 29934 39284 29986
rect 39228 29932 39284 29934
rect 39452 29596 39508 29652
rect 39116 29260 39172 29316
rect 43036 31836 43092 31892
rect 43260 29426 43316 29428
rect 43260 29374 43262 29426
rect 43262 29374 43314 29426
rect 43314 29374 43316 29426
rect 43260 29372 43316 29374
rect 39564 29260 39620 29316
rect 40236 29314 40292 29316
rect 40236 29262 40238 29314
rect 40238 29262 40290 29314
rect 40290 29262 40292 29314
rect 40236 29260 40292 29262
rect 38780 28364 38836 28420
rect 39788 28364 39844 28420
rect 39788 27804 39844 27860
rect 37324 24892 37380 24948
rect 37884 25228 37940 25284
rect 39228 27074 39284 27076
rect 39228 27022 39230 27074
rect 39230 27022 39282 27074
rect 39282 27022 39284 27074
rect 39228 27020 39284 27022
rect 42588 28028 42644 28084
rect 41356 27916 41412 27972
rect 40796 27858 40852 27860
rect 40796 27806 40798 27858
rect 40798 27806 40850 27858
rect 40850 27806 40852 27858
rect 40796 27804 40852 27806
rect 39228 26236 39284 26292
rect 38892 24946 38948 24948
rect 38892 24894 38894 24946
rect 38894 24894 38946 24946
rect 38946 24894 38948 24946
rect 38892 24892 38948 24894
rect 41468 27132 41524 27188
rect 42588 27186 42644 27188
rect 42588 27134 42590 27186
rect 42590 27134 42642 27186
rect 42642 27134 42644 27186
rect 42588 27132 42644 27134
rect 42364 27020 42420 27076
rect 41356 24834 41412 24836
rect 41356 24782 41358 24834
rect 41358 24782 41410 24834
rect 41410 24782 41412 24834
rect 41356 24780 41412 24782
rect 37212 23324 37268 23380
rect 37436 22258 37492 22260
rect 37436 22206 37438 22258
rect 37438 22206 37490 22258
rect 37490 22206 37492 22258
rect 37436 22204 37492 22206
rect 37996 24556 38052 24612
rect 38444 23324 38500 23380
rect 38332 23042 38388 23044
rect 38332 22990 38334 23042
rect 38334 22990 38386 23042
rect 38386 22990 38388 23042
rect 38332 22988 38388 22990
rect 37772 22482 37828 22484
rect 37772 22430 37774 22482
rect 37774 22430 37826 22482
rect 37826 22430 37828 22482
rect 37772 22428 37828 22430
rect 38892 23154 38948 23156
rect 38892 23102 38894 23154
rect 38894 23102 38946 23154
rect 38946 23102 38948 23154
rect 38892 23100 38948 23102
rect 37324 21868 37380 21924
rect 37436 19852 37492 19908
rect 37660 19740 37716 19796
rect 37100 18396 37156 18452
rect 36988 17836 37044 17892
rect 36988 17164 37044 17220
rect 36764 16882 36820 16884
rect 36764 16830 36766 16882
rect 36766 16830 36818 16882
rect 36818 16830 36820 16882
rect 36764 16828 36820 16830
rect 37212 18844 37268 18900
rect 38556 21980 38612 22036
rect 38556 21532 38612 21588
rect 38108 20972 38164 21028
rect 38668 20972 38724 21028
rect 37884 20076 37940 20132
rect 38332 19740 38388 19796
rect 37212 17388 37268 17444
rect 37212 16828 37268 16884
rect 36876 12348 36932 12404
rect 36652 11564 36708 11620
rect 36988 11788 37044 11844
rect 36092 11452 36148 11508
rect 35980 10610 36036 10612
rect 35980 10558 35982 10610
rect 35982 10558 36034 10610
rect 36034 10558 36036 10610
rect 35980 10556 36036 10558
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35868 9938 35924 9940
rect 35868 9886 35870 9938
rect 35870 9886 35922 9938
rect 35922 9886 35924 9938
rect 35868 9884 35924 9886
rect 34860 7644 34916 7700
rect 34300 5010 34356 5012
rect 34300 4958 34302 5010
rect 34302 4958 34354 5010
rect 34354 4958 34356 5010
rect 34300 4956 34356 4958
rect 34076 4562 34132 4564
rect 34076 4510 34078 4562
rect 34078 4510 34130 4562
rect 34130 4510 34132 4562
rect 34076 4508 34132 4510
rect 34524 4450 34580 4452
rect 34524 4398 34526 4450
rect 34526 4398 34578 4450
rect 34578 4398 34580 4450
rect 34524 4396 34580 4398
rect 34300 4338 34356 4340
rect 34300 4286 34302 4338
rect 34302 4286 34354 4338
rect 34354 4286 34356 4338
rect 34300 4284 34356 4286
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35308 8370 35364 8372
rect 35308 8318 35310 8370
rect 35310 8318 35362 8370
rect 35362 8318 35364 8370
rect 35308 8316 35364 8318
rect 36092 9212 36148 9268
rect 36764 9266 36820 9268
rect 36764 9214 36766 9266
rect 36766 9214 36818 9266
rect 36818 9214 36820 9266
rect 36764 9212 36820 9214
rect 36092 8146 36148 8148
rect 36092 8094 36094 8146
rect 36094 8094 36146 8146
rect 36146 8094 36148 8146
rect 36092 8092 36148 8094
rect 35532 7980 35588 8036
rect 36092 7698 36148 7700
rect 36092 7646 36094 7698
rect 36094 7646 36146 7698
rect 36146 7646 36148 7698
rect 36092 7644 36148 7646
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35644 6748 35700 6804
rect 35196 6300 35252 6356
rect 35868 6636 35924 6692
rect 37772 18450 37828 18452
rect 37772 18398 37774 18450
rect 37774 18398 37826 18450
rect 37826 18398 37828 18450
rect 37772 18396 37828 18398
rect 38332 19234 38388 19236
rect 38332 19182 38334 19234
rect 38334 19182 38386 19234
rect 38386 19182 38388 19234
rect 38332 19180 38388 19182
rect 38556 19292 38612 19348
rect 38556 18508 38612 18564
rect 38444 18396 38500 18452
rect 38556 18338 38612 18340
rect 38556 18286 38558 18338
rect 38558 18286 38610 18338
rect 38610 18286 38612 18338
rect 38556 18284 38612 18286
rect 38444 17836 38500 17892
rect 38332 17388 38388 17444
rect 37660 17164 37716 17220
rect 37660 16994 37716 16996
rect 37660 16942 37662 16994
rect 37662 16942 37714 16994
rect 37714 16942 37716 16994
rect 37660 16940 37716 16942
rect 37436 16156 37492 16212
rect 38220 15874 38276 15876
rect 38220 15822 38222 15874
rect 38222 15822 38274 15874
rect 38274 15822 38276 15874
rect 38220 15820 38276 15822
rect 37436 15314 37492 15316
rect 37436 15262 37438 15314
rect 37438 15262 37490 15314
rect 37490 15262 37492 15314
rect 37436 15260 37492 15262
rect 38220 15260 38276 15316
rect 39116 23042 39172 23044
rect 39116 22990 39118 23042
rect 39118 22990 39170 23042
rect 39170 22990 39172 23042
rect 39116 22988 39172 22990
rect 40572 24556 40628 24612
rect 39340 21196 39396 21252
rect 37772 13858 37828 13860
rect 37772 13806 37774 13858
rect 37774 13806 37826 13858
rect 37826 13806 37828 13858
rect 37772 13804 37828 13806
rect 37996 13692 38052 13748
rect 37324 11564 37380 11620
rect 38556 14924 38612 14980
rect 38556 14642 38612 14644
rect 38556 14590 38558 14642
rect 38558 14590 38610 14642
rect 38610 14590 38612 14642
rect 38556 14588 38612 14590
rect 38668 14418 38724 14420
rect 38668 14366 38670 14418
rect 38670 14366 38722 14418
rect 38722 14366 38724 14418
rect 38668 14364 38724 14366
rect 38668 13692 38724 13748
rect 39340 20018 39396 20020
rect 39340 19966 39342 20018
rect 39342 19966 39394 20018
rect 39394 19966 39396 20018
rect 39340 19964 39396 19966
rect 40236 20748 40292 20804
rect 40012 19852 40068 19908
rect 40124 20076 40180 20132
rect 40460 19964 40516 20020
rect 39452 18844 39508 18900
rect 40124 18844 40180 18900
rect 39228 18450 39284 18452
rect 39228 18398 39230 18450
rect 39230 18398 39282 18450
rect 39282 18398 39284 18450
rect 39228 18396 39284 18398
rect 39340 18284 39396 18340
rect 40124 18338 40180 18340
rect 40124 18286 40126 18338
rect 40126 18286 40178 18338
rect 40178 18286 40180 18338
rect 40124 18284 40180 18286
rect 41692 24610 41748 24612
rect 41692 24558 41694 24610
rect 41694 24558 41746 24610
rect 41746 24558 41748 24610
rect 41692 24556 41748 24558
rect 42252 26290 42308 26292
rect 42252 26238 42254 26290
rect 42254 26238 42306 26290
rect 42306 26238 42308 26290
rect 42252 26236 42308 26238
rect 43596 33180 43652 33236
rect 43708 32956 43764 33012
rect 43932 32674 43988 32676
rect 43932 32622 43934 32674
rect 43934 32622 43986 32674
rect 43986 32622 43988 32674
rect 43932 32620 43988 32622
rect 43708 31836 43764 31892
rect 44268 36988 44324 37044
rect 44156 36652 44212 36708
rect 44492 37266 44548 37268
rect 44492 37214 44494 37266
rect 44494 37214 44546 37266
rect 44546 37214 44548 37266
rect 44492 37212 44548 37214
rect 46284 40402 46340 40404
rect 46284 40350 46286 40402
rect 46286 40350 46338 40402
rect 46338 40350 46340 40402
rect 46284 40348 46340 40350
rect 46060 39564 46116 39620
rect 45612 38946 45668 38948
rect 45612 38894 45614 38946
rect 45614 38894 45666 38946
rect 45666 38894 45668 38946
rect 45612 38892 45668 38894
rect 45948 39004 46004 39060
rect 45164 38834 45220 38836
rect 45164 38782 45166 38834
rect 45166 38782 45218 38834
rect 45218 38782 45220 38834
rect 45164 38780 45220 38782
rect 46284 39340 46340 39396
rect 46396 38834 46452 38836
rect 46396 38782 46398 38834
rect 46398 38782 46450 38834
rect 46450 38782 46452 38834
rect 46396 38780 46452 38782
rect 47516 42082 47572 42084
rect 47516 42030 47518 42082
rect 47518 42030 47570 42082
rect 47570 42030 47572 42082
rect 47516 42028 47572 42030
rect 47292 41970 47348 41972
rect 47292 41918 47294 41970
rect 47294 41918 47346 41970
rect 47346 41918 47348 41970
rect 47292 41916 47348 41918
rect 46732 41580 46788 41636
rect 46620 41298 46676 41300
rect 46620 41246 46622 41298
rect 46622 41246 46674 41298
rect 46674 41246 46676 41298
rect 46620 41244 46676 41246
rect 46732 40908 46788 40964
rect 47068 41356 47124 41412
rect 47292 41692 47348 41748
rect 48412 48300 48468 48356
rect 47740 48130 47796 48132
rect 47740 48078 47742 48130
rect 47742 48078 47794 48130
rect 47794 48078 47796 48130
rect 47740 48076 47796 48078
rect 47964 48188 48020 48244
rect 47852 48018 47908 48020
rect 47852 47966 47854 48018
rect 47854 47966 47906 48018
rect 47906 47966 47908 48018
rect 47852 47964 47908 47966
rect 48076 45948 48132 46004
rect 48412 45276 48468 45332
rect 47740 45218 47796 45220
rect 47740 45166 47742 45218
rect 47742 45166 47794 45218
rect 47794 45166 47796 45218
rect 47740 45164 47796 45166
rect 48412 43708 48468 43764
rect 47740 43484 47796 43540
rect 47852 41970 47908 41972
rect 47852 41918 47854 41970
rect 47854 41918 47906 41970
rect 47906 41918 47908 41970
rect 47852 41916 47908 41918
rect 47628 41132 47684 41188
rect 46620 39340 46676 39396
rect 46844 39394 46900 39396
rect 46844 39342 46846 39394
rect 46846 39342 46898 39394
rect 46898 39342 46900 39394
rect 46844 39340 46900 39342
rect 45052 37436 45108 37492
rect 44940 36988 44996 37044
rect 44716 36652 44772 36708
rect 44828 35420 44884 35476
rect 44940 36316 44996 36372
rect 45724 37266 45780 37268
rect 45724 37214 45726 37266
rect 45726 37214 45778 37266
rect 45778 37214 45780 37266
rect 45724 37212 45780 37214
rect 45948 37266 46004 37268
rect 45948 37214 45950 37266
rect 45950 37214 46002 37266
rect 46002 37214 46004 37266
rect 45948 37212 46004 37214
rect 45388 36988 45444 37044
rect 45276 36428 45332 36484
rect 45724 35532 45780 35588
rect 45164 34748 45220 34804
rect 44604 33516 44660 33572
rect 45388 33628 45444 33684
rect 45276 33346 45332 33348
rect 45276 33294 45278 33346
rect 45278 33294 45330 33346
rect 45330 33294 45332 33346
rect 45276 33292 45332 33294
rect 44044 31724 44100 31780
rect 44156 31836 44212 31892
rect 45612 33180 45668 33236
rect 45388 31218 45444 31220
rect 45388 31166 45390 31218
rect 45390 31166 45442 31218
rect 45442 31166 45444 31218
rect 45388 31164 45444 31166
rect 44268 30098 44324 30100
rect 44268 30046 44270 30098
rect 44270 30046 44322 30098
rect 44322 30046 44324 30098
rect 44268 30044 44324 30046
rect 45612 30098 45668 30100
rect 45612 30046 45614 30098
rect 45614 30046 45666 30098
rect 45666 30046 45668 30098
rect 45612 30044 45668 30046
rect 46060 36652 46116 36708
rect 46060 36482 46116 36484
rect 46060 36430 46062 36482
rect 46062 36430 46114 36482
rect 46114 36430 46116 36482
rect 46060 36428 46116 36430
rect 45948 33292 46004 33348
rect 47292 40236 47348 40292
rect 46956 37212 47012 37268
rect 47180 36652 47236 36708
rect 47292 36370 47348 36372
rect 47292 36318 47294 36370
rect 47294 36318 47346 36370
rect 47346 36318 47348 36370
rect 47292 36316 47348 36318
rect 46732 35586 46788 35588
rect 46732 35534 46734 35586
rect 46734 35534 46786 35586
rect 46786 35534 46788 35586
rect 46732 35532 46788 35534
rect 47068 34972 47124 35028
rect 46844 34914 46900 34916
rect 46844 34862 46846 34914
rect 46846 34862 46898 34914
rect 46898 34862 46900 34914
rect 46844 34860 46900 34862
rect 46508 34354 46564 34356
rect 46508 34302 46510 34354
rect 46510 34302 46562 34354
rect 46562 34302 46564 34354
rect 46508 34300 46564 34302
rect 47404 35868 47460 35924
rect 47516 35084 47572 35140
rect 48188 42140 48244 42196
rect 48412 42028 48468 42084
rect 48076 41298 48132 41300
rect 48076 41246 48078 41298
rect 48078 41246 48130 41298
rect 48130 41246 48132 41298
rect 48076 41244 48132 41246
rect 47852 41020 47908 41076
rect 48188 40962 48244 40964
rect 48188 40910 48190 40962
rect 48190 40910 48242 40962
rect 48242 40910 48244 40962
rect 48188 40908 48244 40910
rect 48412 39618 48468 39620
rect 48412 39566 48414 39618
rect 48414 39566 48466 39618
rect 48466 39566 48468 39618
rect 48412 39564 48468 39566
rect 47852 39058 47908 39060
rect 47852 39006 47854 39058
rect 47854 39006 47906 39058
rect 47906 39006 47908 39058
rect 47852 39004 47908 39006
rect 48860 50428 48916 50484
rect 48972 48242 49028 48244
rect 48972 48190 48974 48242
rect 48974 48190 49026 48242
rect 49026 48190 49028 48242
rect 48972 48188 49028 48190
rect 48860 47964 48916 48020
rect 48748 47068 48804 47124
rect 48972 47404 49028 47460
rect 49084 46786 49140 46788
rect 49084 46734 49086 46786
rect 49086 46734 49138 46786
rect 49138 46734 49140 46786
rect 49084 46732 49140 46734
rect 49868 54290 49924 54292
rect 49868 54238 49870 54290
rect 49870 54238 49922 54290
rect 49922 54238 49924 54290
rect 49868 54236 49924 54238
rect 50092 53564 50148 53620
rect 50092 53004 50148 53060
rect 50652 54514 50708 54516
rect 50652 54462 50654 54514
rect 50654 54462 50706 54514
rect 50706 54462 50708 54514
rect 50652 54460 50708 54462
rect 54012 56082 54068 56084
rect 54012 56030 54014 56082
rect 54014 56030 54066 56082
rect 54066 56030 54068 56082
rect 54012 56028 54068 56030
rect 51436 54684 51492 54740
rect 51884 54684 51940 54740
rect 50876 54348 50932 54404
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 51100 53676 51156 53732
rect 52780 53676 52836 53732
rect 50204 52220 50260 52276
rect 50428 52108 50484 52164
rect 50988 52162 51044 52164
rect 50988 52110 50990 52162
rect 50990 52110 51042 52162
rect 51042 52110 51044 52162
rect 50988 52108 51044 52110
rect 50316 51996 50372 52052
rect 51548 53058 51604 53060
rect 51548 53006 51550 53058
rect 51550 53006 51602 53058
rect 51602 53006 51604 53058
rect 51548 53004 51604 53006
rect 51212 52050 51268 52052
rect 51212 51998 51214 52050
rect 51214 51998 51266 52050
rect 51266 51998 51268 52050
rect 51212 51996 51268 51998
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 49644 50706 49700 50708
rect 49644 50654 49646 50706
rect 49646 50654 49698 50706
rect 49698 50654 49700 50706
rect 49644 50652 49700 50654
rect 50652 50652 50708 50708
rect 50092 50594 50148 50596
rect 50092 50542 50094 50594
rect 50094 50542 50146 50594
rect 50146 50542 50148 50594
rect 50092 50540 50148 50542
rect 51212 50652 51268 50708
rect 54572 54514 54628 54516
rect 54572 54462 54574 54514
rect 54574 54462 54626 54514
rect 54626 54462 54628 54514
rect 54572 54460 54628 54462
rect 53228 54348 53284 54404
rect 53900 53676 53956 53732
rect 55580 53730 55636 53732
rect 55580 53678 55582 53730
rect 55582 53678 55634 53730
rect 55634 53678 55636 53730
rect 55580 53676 55636 53678
rect 57260 53116 57316 53172
rect 51996 50652 52052 50708
rect 52332 50652 52388 50708
rect 49420 50428 49476 50484
rect 50204 50482 50260 50484
rect 50204 50430 50206 50482
rect 50206 50430 50258 50482
rect 50258 50430 50260 50482
rect 50204 50428 50260 50430
rect 50764 50482 50820 50484
rect 50764 50430 50766 50482
rect 50766 50430 50818 50482
rect 50818 50430 50820 50482
rect 50764 50428 50820 50430
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 52668 50706 52724 50708
rect 52668 50654 52670 50706
rect 52670 50654 52722 50706
rect 52722 50654 52724 50706
rect 52668 50652 52724 50654
rect 52892 50316 52948 50372
rect 51772 49810 51828 49812
rect 51772 49758 51774 49810
rect 51774 49758 51826 49810
rect 51826 49758 51828 49810
rect 51772 49756 51828 49758
rect 53004 49756 53060 49812
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 49420 48354 49476 48356
rect 49420 48302 49422 48354
rect 49422 48302 49474 48354
rect 49474 48302 49476 48354
rect 49420 48300 49476 48302
rect 53116 49138 53172 49140
rect 53116 49086 53118 49138
rect 53118 49086 53170 49138
rect 53170 49086 53172 49138
rect 53116 49084 53172 49086
rect 54348 50316 54404 50372
rect 53900 49810 53956 49812
rect 53900 49758 53902 49810
rect 53902 49758 53954 49810
rect 53954 49758 53956 49810
rect 53900 49756 53956 49758
rect 54236 49868 54292 49924
rect 53900 49138 53956 49140
rect 53900 49086 53902 49138
rect 53902 49086 53954 49138
rect 53954 49086 53956 49138
rect 53900 49084 53956 49086
rect 53676 48972 53732 49028
rect 51996 48802 52052 48804
rect 51996 48750 51998 48802
rect 51998 48750 52050 48802
rect 52050 48750 52052 48802
rect 51996 48748 52052 48750
rect 52780 48802 52836 48804
rect 52780 48750 52782 48802
rect 52782 48750 52834 48802
rect 52834 48750 52836 48802
rect 52780 48748 52836 48750
rect 49532 47628 49588 47684
rect 48748 45948 48804 46004
rect 48748 45778 48804 45780
rect 48748 45726 48750 45778
rect 48750 45726 48802 45778
rect 48802 45726 48804 45778
rect 48748 45724 48804 45726
rect 48748 45106 48804 45108
rect 48748 45054 48750 45106
rect 48750 45054 48802 45106
rect 48802 45054 48804 45106
rect 48748 45052 48804 45054
rect 49196 45724 49252 45780
rect 48972 45218 49028 45220
rect 48972 45166 48974 45218
rect 48974 45166 49026 45218
rect 49026 45166 49028 45218
rect 48972 45164 49028 45166
rect 49084 43538 49140 43540
rect 49084 43486 49086 43538
rect 49086 43486 49138 43538
rect 49138 43486 49140 43538
rect 49084 43484 49140 43486
rect 48860 42530 48916 42532
rect 48860 42478 48862 42530
rect 48862 42478 48914 42530
rect 48914 42478 48916 42530
rect 48860 42476 48916 42478
rect 49308 45276 49364 45332
rect 50204 47458 50260 47460
rect 50204 47406 50206 47458
rect 50206 47406 50258 47458
rect 50258 47406 50260 47458
rect 50204 47404 50260 47406
rect 49756 47068 49812 47124
rect 50428 48188 50484 48244
rect 50316 46786 50372 46788
rect 50316 46734 50318 46786
rect 50318 46734 50370 46786
rect 50370 46734 50372 46786
rect 50316 46732 50372 46734
rect 49644 45778 49700 45780
rect 49644 45726 49646 45778
rect 49646 45726 49698 45778
rect 49698 45726 49700 45778
rect 49644 45724 49700 45726
rect 49980 44994 50036 44996
rect 49980 44942 49982 44994
rect 49982 44942 50034 44994
rect 50034 44942 50036 44994
rect 49980 44940 50036 44942
rect 49420 42924 49476 42980
rect 50764 47628 50820 47684
rect 52108 47404 52164 47460
rect 52444 48242 52500 48244
rect 52444 48190 52446 48242
rect 52446 48190 52498 48242
rect 52498 48190 52500 48242
rect 52444 48188 52500 48190
rect 51772 47234 51828 47236
rect 51772 47182 51774 47234
rect 51774 47182 51826 47234
rect 51826 47182 51828 47234
rect 51772 47180 51828 47182
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 50988 47068 51044 47124
rect 52220 47180 52276 47236
rect 51996 47068 52052 47124
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 50316 45164 50372 45220
rect 50764 44994 50820 44996
rect 50764 44942 50766 44994
rect 50766 44942 50818 44994
rect 50818 44942 50820 44994
rect 50764 44940 50820 44942
rect 50652 44380 50708 44436
rect 50988 44380 51044 44436
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 50092 43708 50148 43764
rect 52332 46674 52388 46676
rect 52332 46622 52334 46674
rect 52334 46622 52386 46674
rect 52386 46622 52388 46674
rect 52332 46620 52388 46622
rect 52668 47964 52724 48020
rect 52668 47068 52724 47124
rect 53228 48188 53284 48244
rect 53004 48018 53060 48020
rect 53004 47966 53006 48018
rect 53006 47966 53058 48018
rect 53058 47966 53060 48018
rect 53004 47964 53060 47966
rect 52892 47404 52948 47460
rect 53564 46674 53620 46676
rect 53564 46622 53566 46674
rect 53566 46622 53618 46674
rect 53618 46622 53620 46674
rect 53564 46620 53620 46622
rect 54236 49026 54292 49028
rect 54236 48974 54238 49026
rect 54238 48974 54290 49026
rect 54290 48974 54292 49026
rect 54236 48972 54292 48974
rect 54908 49922 54964 49924
rect 54908 49870 54910 49922
rect 54910 49870 54962 49922
rect 54962 49870 54964 49922
rect 54908 49868 54964 49870
rect 57820 50316 57876 50372
rect 57932 49756 57988 49812
rect 58156 47068 58212 47124
rect 53116 44268 53172 44324
rect 51212 43596 51268 43652
rect 49868 42812 49924 42868
rect 49420 42754 49476 42756
rect 49420 42702 49422 42754
rect 49422 42702 49474 42754
rect 49474 42702 49476 42754
rect 49420 42700 49476 42702
rect 48636 41186 48692 41188
rect 48636 41134 48638 41186
rect 48638 41134 48690 41186
rect 48690 41134 48692 41186
rect 48636 41132 48692 41134
rect 49084 42194 49140 42196
rect 49084 42142 49086 42194
rect 49086 42142 49138 42194
rect 49138 42142 49140 42194
rect 49084 42140 49140 42142
rect 49308 42082 49364 42084
rect 49308 42030 49310 42082
rect 49310 42030 49362 42082
rect 49362 42030 49364 42082
rect 49308 42028 49364 42030
rect 48972 41916 49028 41972
rect 49196 41970 49252 41972
rect 49196 41918 49198 41970
rect 49198 41918 49250 41970
rect 49250 41918 49252 41970
rect 49196 41916 49252 41918
rect 49980 42924 50036 42980
rect 51212 42866 51268 42868
rect 51212 42814 51214 42866
rect 51214 42814 51266 42866
rect 51266 42814 51268 42866
rect 51212 42812 51268 42814
rect 50092 42700 50148 42756
rect 49084 41298 49140 41300
rect 49084 41246 49086 41298
rect 49086 41246 49138 41298
rect 49138 41246 49140 41298
rect 49084 41244 49140 41246
rect 48748 41020 48804 41076
rect 48636 39340 48692 39396
rect 47628 34972 47684 35028
rect 49084 39842 49140 39844
rect 49084 39790 49086 39842
rect 49086 39790 49138 39842
rect 49138 39790 49140 39842
rect 49084 39788 49140 39790
rect 48972 39506 49028 39508
rect 48972 39454 48974 39506
rect 48974 39454 49026 39506
rect 49026 39454 49028 39506
rect 48972 39452 49028 39454
rect 48972 39004 49028 39060
rect 49420 40514 49476 40516
rect 49420 40462 49422 40514
rect 49422 40462 49474 40514
rect 49474 40462 49476 40514
rect 49420 40460 49476 40462
rect 49532 39788 49588 39844
rect 49980 41244 50036 41300
rect 49756 39564 49812 39620
rect 49644 39506 49700 39508
rect 49644 39454 49646 39506
rect 49646 39454 49698 39506
rect 49698 39454 49700 39506
rect 49644 39452 49700 39454
rect 49868 39340 49924 39396
rect 50092 39452 50148 39508
rect 49308 39004 49364 39060
rect 49644 39058 49700 39060
rect 49644 39006 49646 39058
rect 49646 39006 49698 39058
rect 49698 39006 49700 39058
rect 49644 39004 49700 39006
rect 50092 38892 50148 38948
rect 48748 38722 48804 38724
rect 48748 38670 48750 38722
rect 48750 38670 48802 38722
rect 48802 38670 48804 38722
rect 48748 38668 48804 38670
rect 46844 34300 46900 34356
rect 46284 33180 46340 33236
rect 47516 33404 47572 33460
rect 47180 33346 47236 33348
rect 47180 33294 47182 33346
rect 47182 33294 47234 33346
rect 47234 33294 47236 33346
rect 47180 33292 47236 33294
rect 47068 33180 47124 33236
rect 46956 32674 47012 32676
rect 46956 32622 46958 32674
rect 46958 32622 47010 32674
rect 47010 32622 47012 32674
rect 46956 32620 47012 32622
rect 47516 32786 47572 32788
rect 47516 32734 47518 32786
rect 47518 32734 47570 32786
rect 47570 32734 47572 32786
rect 47516 32732 47572 32734
rect 47628 32620 47684 32676
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 51772 43596 51828 43652
rect 51660 43538 51716 43540
rect 51660 43486 51662 43538
rect 51662 43486 51714 43538
rect 51714 43486 51716 43538
rect 51660 43484 51716 43486
rect 52220 43596 52276 43652
rect 53900 43650 53956 43652
rect 53900 43598 53902 43650
rect 53902 43598 53954 43650
rect 53954 43598 53956 43650
rect 53900 43596 53956 43598
rect 52332 43484 52388 43540
rect 52892 43484 52948 43540
rect 51772 42700 51828 42756
rect 51548 42476 51604 42532
rect 51884 42140 51940 42196
rect 51212 41970 51268 41972
rect 51212 41918 51214 41970
rect 51214 41918 51266 41970
rect 51266 41918 51268 41970
rect 51212 41916 51268 41918
rect 51436 41916 51492 41972
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 50540 40514 50596 40516
rect 50540 40462 50542 40514
rect 50542 40462 50594 40514
rect 50594 40462 50596 40514
rect 50540 40460 50596 40462
rect 50764 39900 50820 39956
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 50540 38946 50596 38948
rect 50540 38894 50542 38946
rect 50542 38894 50594 38946
rect 50594 38894 50596 38946
rect 50540 38892 50596 38894
rect 50988 40908 51044 40964
rect 52556 42194 52612 42196
rect 52556 42142 52558 42194
rect 52558 42142 52610 42194
rect 52610 42142 52612 42194
rect 52556 42140 52612 42142
rect 52444 41970 52500 41972
rect 52444 41918 52446 41970
rect 52446 41918 52498 41970
rect 52498 41918 52500 41970
rect 52444 41916 52500 41918
rect 51772 41074 51828 41076
rect 51772 41022 51774 41074
rect 51774 41022 51826 41074
rect 51826 41022 51828 41074
rect 51772 41020 51828 41022
rect 53004 42754 53060 42756
rect 53004 42702 53006 42754
rect 53006 42702 53058 42754
rect 53058 42702 53060 42754
rect 53004 42700 53060 42702
rect 54572 44322 54628 44324
rect 54572 44270 54574 44322
rect 54574 44270 54626 44322
rect 54626 44270 54628 44322
rect 54572 44268 54628 44270
rect 54460 43596 54516 43652
rect 53452 42140 53508 42196
rect 57932 44434 57988 44436
rect 57932 44382 57934 44434
rect 57934 44382 57986 44434
rect 57986 44382 57988 44434
rect 57932 44380 57988 44382
rect 54796 43538 54852 43540
rect 54796 43486 54798 43538
rect 54798 43486 54850 43538
rect 54850 43486 54852 43538
rect 54796 43484 54852 43486
rect 55468 43538 55524 43540
rect 55468 43486 55470 43538
rect 55470 43486 55522 43538
rect 55522 43486 55524 43538
rect 55468 43484 55524 43486
rect 56812 43538 56868 43540
rect 56812 43486 56814 43538
rect 56814 43486 56866 43538
rect 56866 43486 56868 43538
rect 56812 43484 56868 43486
rect 57932 43036 57988 43092
rect 53004 41074 53060 41076
rect 53004 41022 53006 41074
rect 53006 41022 53058 41074
rect 53058 41022 53060 41074
rect 53004 41020 53060 41022
rect 54348 41074 54404 41076
rect 54348 41022 54350 41074
rect 54350 41022 54402 41074
rect 54402 41022 54404 41074
rect 54348 41020 54404 41022
rect 51660 40514 51716 40516
rect 51660 40462 51662 40514
rect 51662 40462 51714 40514
rect 51714 40462 51716 40514
rect 51660 40460 51716 40462
rect 53676 40626 53732 40628
rect 53676 40574 53678 40626
rect 53678 40574 53730 40626
rect 53730 40574 53732 40626
rect 53676 40572 53732 40574
rect 54460 40572 54516 40628
rect 55132 41020 55188 41076
rect 55020 40236 55076 40292
rect 51100 39900 51156 39956
rect 50988 39506 51044 39508
rect 50988 39454 50990 39506
rect 50990 39454 51042 39506
rect 51042 39454 51044 39506
rect 50988 39452 51044 39454
rect 51100 39004 51156 39060
rect 53228 39452 53284 39508
rect 53228 39058 53284 39060
rect 53228 39006 53230 39058
rect 53230 39006 53282 39058
rect 53282 39006 53284 39058
rect 53228 39004 53284 39006
rect 51884 38780 51940 38836
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 49756 37378 49812 37380
rect 49756 37326 49758 37378
rect 49758 37326 49810 37378
rect 49810 37326 49812 37378
rect 49756 37324 49812 37326
rect 50092 37266 50148 37268
rect 50092 37214 50094 37266
rect 50094 37214 50146 37266
rect 50146 37214 50148 37266
rect 50092 37212 50148 37214
rect 49868 37154 49924 37156
rect 49868 37102 49870 37154
rect 49870 37102 49922 37154
rect 49922 37102 49924 37154
rect 49868 37100 49924 37102
rect 47852 35868 47908 35924
rect 48076 35810 48132 35812
rect 48076 35758 48078 35810
rect 48078 35758 48130 35810
rect 48130 35758 48132 35810
rect 48076 35756 48132 35758
rect 49084 35698 49140 35700
rect 49084 35646 49086 35698
rect 49086 35646 49138 35698
rect 49138 35646 49140 35698
rect 49084 35644 49140 35646
rect 48860 35420 48916 35476
rect 49532 35756 49588 35812
rect 50652 37490 50708 37492
rect 50652 37438 50654 37490
rect 50654 37438 50706 37490
rect 50706 37438 50708 37490
rect 50652 37436 50708 37438
rect 50540 37212 50596 37268
rect 53116 38834 53172 38836
rect 53116 38782 53118 38834
rect 53118 38782 53170 38834
rect 53170 38782 53172 38834
rect 53116 38780 53172 38782
rect 51660 37378 51716 37380
rect 51660 37326 51662 37378
rect 51662 37326 51714 37378
rect 51714 37326 51716 37378
rect 51660 37324 51716 37326
rect 52892 37266 52948 37268
rect 52892 37214 52894 37266
rect 52894 37214 52946 37266
rect 52946 37214 52948 37266
rect 52892 37212 52948 37214
rect 51436 37100 51492 37156
rect 53004 36316 53060 36372
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 49308 35084 49364 35140
rect 50428 35084 50484 35140
rect 48076 34972 48132 35028
rect 50316 35026 50372 35028
rect 50316 34974 50318 35026
rect 50318 34974 50370 35026
rect 50370 34974 50372 35026
rect 50316 34972 50372 34974
rect 48748 34914 48804 34916
rect 48748 34862 48750 34914
rect 48750 34862 48802 34914
rect 48802 34862 48804 34914
rect 48748 34860 48804 34862
rect 49196 34636 49252 34692
rect 51996 34748 52052 34804
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 50876 34354 50932 34356
rect 50876 34302 50878 34354
rect 50878 34302 50930 34354
rect 50930 34302 50932 34354
rect 50876 34300 50932 34302
rect 51436 34300 51492 34356
rect 50652 34242 50708 34244
rect 50652 34190 50654 34242
rect 50654 34190 50706 34242
rect 50706 34190 50708 34242
rect 50652 34188 50708 34190
rect 50092 34130 50148 34132
rect 50092 34078 50094 34130
rect 50094 34078 50146 34130
rect 50146 34078 50148 34130
rect 50092 34076 50148 34078
rect 50764 34130 50820 34132
rect 50764 34078 50766 34130
rect 50766 34078 50818 34130
rect 50818 34078 50820 34130
rect 50764 34076 50820 34078
rect 48636 33346 48692 33348
rect 48636 33294 48638 33346
rect 48638 33294 48690 33346
rect 48690 33294 48692 33346
rect 48636 33292 48692 33294
rect 49532 33346 49588 33348
rect 49532 33294 49534 33346
rect 49534 33294 49586 33346
rect 49586 33294 49588 33346
rect 49532 33292 49588 33294
rect 48188 33234 48244 33236
rect 48188 33182 48190 33234
rect 48190 33182 48242 33234
rect 48242 33182 48244 33234
rect 48188 33180 48244 33182
rect 48076 32786 48132 32788
rect 48076 32734 48078 32786
rect 48078 32734 48130 32786
rect 48130 32734 48132 32786
rect 48076 32732 48132 32734
rect 48524 33234 48580 33236
rect 48524 33182 48526 33234
rect 48526 33182 48578 33234
rect 48578 33182 48580 33234
rect 48524 33180 48580 33182
rect 48188 31948 48244 32004
rect 48860 32002 48916 32004
rect 48860 31950 48862 32002
rect 48862 31950 48914 32002
rect 48914 31950 48916 32002
rect 48860 31948 48916 31950
rect 49196 32732 49252 32788
rect 52780 35196 52836 35252
rect 53228 35698 53284 35700
rect 53228 35646 53230 35698
rect 53230 35646 53282 35698
rect 53282 35646 53284 35698
rect 53228 35644 53284 35646
rect 53452 38050 53508 38052
rect 53452 37998 53454 38050
rect 53454 37998 53506 38050
rect 53506 37998 53508 38050
rect 53452 37996 53508 37998
rect 54124 39004 54180 39060
rect 53900 37436 53956 37492
rect 54012 38780 54068 38836
rect 54572 39004 54628 39060
rect 55244 40348 55300 40404
rect 56924 40402 56980 40404
rect 56924 40350 56926 40402
rect 56926 40350 56978 40402
rect 56978 40350 56980 40402
rect 56924 40348 56980 40350
rect 57932 40348 57988 40404
rect 56812 40290 56868 40292
rect 56812 40238 56814 40290
rect 56814 40238 56866 40290
rect 56866 40238 56868 40290
rect 56812 40236 56868 40238
rect 54796 37996 54852 38052
rect 54348 36370 54404 36372
rect 54348 36318 54350 36370
rect 54350 36318 54402 36370
rect 54402 36318 54404 36370
rect 54348 36316 54404 36318
rect 53788 35644 53844 35700
rect 53340 35196 53396 35252
rect 52780 34802 52836 34804
rect 52780 34750 52782 34802
rect 52782 34750 52834 34802
rect 52834 34750 52836 34802
rect 52780 34748 52836 34750
rect 52892 34690 52948 34692
rect 52892 34638 52894 34690
rect 52894 34638 52946 34690
rect 52946 34638 52948 34690
rect 52892 34636 52948 34638
rect 52444 34188 52500 34244
rect 50764 33458 50820 33460
rect 50764 33406 50766 33458
rect 50766 33406 50818 33458
rect 50818 33406 50820 33458
rect 50764 33404 50820 33406
rect 50204 33292 50260 33348
rect 50876 33292 50932 33348
rect 50092 33068 50148 33124
rect 49644 32732 49700 32788
rect 53004 34300 53060 34356
rect 54236 35698 54292 35700
rect 54236 35646 54238 35698
rect 54238 35646 54290 35698
rect 54290 35646 54292 35698
rect 54236 35644 54292 35646
rect 54236 35196 54292 35252
rect 55356 36204 55412 36260
rect 54684 35644 54740 35700
rect 54460 34748 54516 34804
rect 55356 34972 55412 35028
rect 56588 36258 56644 36260
rect 56588 36206 56590 36258
rect 56590 36206 56642 36258
rect 56642 36206 56644 36258
rect 56588 36204 56644 36206
rect 57932 37660 57988 37716
rect 57708 35644 57764 35700
rect 55804 35420 55860 35476
rect 55804 34802 55860 34804
rect 55804 34750 55806 34802
rect 55806 34750 55858 34802
rect 55858 34750 55860 34802
rect 55804 34748 55860 34750
rect 51884 33292 51940 33348
rect 53004 33346 53060 33348
rect 53004 33294 53006 33346
rect 53006 33294 53058 33346
rect 53058 33294 53060 33346
rect 53004 33292 53060 33294
rect 54348 33292 54404 33348
rect 51324 33234 51380 33236
rect 51324 33182 51326 33234
rect 51326 33182 51378 33234
rect 51378 33182 51380 33234
rect 51324 33180 51380 33182
rect 55580 33346 55636 33348
rect 55580 33294 55582 33346
rect 55582 33294 55634 33346
rect 55634 33294 55636 33346
rect 55580 33292 55636 33294
rect 51436 33122 51492 33124
rect 51436 33070 51438 33122
rect 51438 33070 51490 33122
rect 51490 33070 51492 33122
rect 51436 33068 51492 33070
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 57932 32956 57988 33012
rect 50764 32900 50820 32902
rect 49532 32508 49588 32564
rect 49868 32562 49924 32564
rect 49868 32510 49870 32562
rect 49870 32510 49922 32562
rect 49922 32510 49924 32562
rect 49868 32508 49924 32510
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 57820 31106 57876 31108
rect 57820 31054 57822 31106
rect 57822 31054 57874 31106
rect 57874 31054 57876 31106
rect 57820 31052 57876 31054
rect 58156 30268 58212 30324
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 43932 29372 43988 29428
rect 43932 28082 43988 28084
rect 43932 28030 43934 28082
rect 43934 28030 43986 28082
rect 43986 28030 43988 28082
rect 43932 28028 43988 28030
rect 45164 28028 45220 28084
rect 44492 27634 44548 27636
rect 44492 27582 44494 27634
rect 44494 27582 44546 27634
rect 44546 27582 44548 27634
rect 44492 27580 44548 27582
rect 43484 27074 43540 27076
rect 43484 27022 43486 27074
rect 43486 27022 43538 27074
rect 43538 27022 43540 27074
rect 43484 27020 43540 27022
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 58156 28252 58212 28308
rect 50764 28196 50820 28198
rect 45612 28028 45668 28084
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 43484 26012 43540 26068
rect 43372 25452 43428 25508
rect 42700 25228 42756 25284
rect 41132 23772 41188 23828
rect 40908 23378 40964 23380
rect 40908 23326 40910 23378
rect 40910 23326 40962 23378
rect 40962 23326 40964 23378
rect 40908 23324 40964 23326
rect 41804 23660 41860 23716
rect 41692 23548 41748 23604
rect 40796 22092 40852 22148
rect 40684 19458 40740 19460
rect 40684 19406 40686 19458
rect 40686 19406 40738 19458
rect 40738 19406 40740 19458
rect 40684 19404 40740 19406
rect 41132 21196 41188 21252
rect 41132 20524 41188 20580
rect 40908 20300 40964 20356
rect 42812 25116 42868 25172
rect 45948 26066 46004 26068
rect 45948 26014 45950 26066
rect 45950 26014 46002 26066
rect 46002 26014 46004 26066
rect 45948 26012 46004 26014
rect 43932 25506 43988 25508
rect 43932 25454 43934 25506
rect 43934 25454 43986 25506
rect 43986 25454 43988 25506
rect 43932 25452 43988 25454
rect 43484 25228 43540 25284
rect 44828 25116 44884 25172
rect 42140 23772 42196 23828
rect 42252 23884 42308 23940
rect 42476 23714 42532 23716
rect 42476 23662 42478 23714
rect 42478 23662 42530 23714
rect 42530 23662 42532 23714
rect 42476 23660 42532 23662
rect 42364 23548 42420 23604
rect 42700 23548 42756 23604
rect 41916 22204 41972 22260
rect 41356 20860 41412 20916
rect 41580 21586 41636 21588
rect 41580 21534 41582 21586
rect 41582 21534 41634 21586
rect 41634 21534 41636 21586
rect 41580 21532 41636 21534
rect 41580 20802 41636 20804
rect 41580 20750 41582 20802
rect 41582 20750 41634 20802
rect 41634 20750 41636 20802
rect 41580 20748 41636 20750
rect 41468 20636 41524 20692
rect 41580 20524 41636 20580
rect 40796 18956 40852 19012
rect 41692 19964 41748 20020
rect 41692 19404 41748 19460
rect 41580 18956 41636 19012
rect 39116 17442 39172 17444
rect 39116 17390 39118 17442
rect 39118 17390 39170 17442
rect 39170 17390 39172 17442
rect 39116 17388 39172 17390
rect 39004 14476 39060 14532
rect 39900 15820 39956 15876
rect 40124 16044 40180 16100
rect 39228 15036 39284 15092
rect 39788 15036 39844 15092
rect 39452 14530 39508 14532
rect 39452 14478 39454 14530
rect 39454 14478 39506 14530
rect 39506 14478 39508 14530
rect 39452 14476 39508 14478
rect 39116 14364 39172 14420
rect 38892 13804 38948 13860
rect 39340 13858 39396 13860
rect 39340 13806 39342 13858
rect 39342 13806 39394 13858
rect 39394 13806 39396 13858
rect 39340 13804 39396 13806
rect 37212 10556 37268 10612
rect 40236 15090 40292 15092
rect 40236 15038 40238 15090
rect 40238 15038 40290 15090
rect 40290 15038 40292 15090
rect 40236 15036 40292 15038
rect 38780 11676 38836 11732
rect 37548 10444 37604 10500
rect 37212 9884 37268 9940
rect 37100 9212 37156 9268
rect 36204 5906 36260 5908
rect 36204 5854 36206 5906
rect 36206 5854 36258 5906
rect 36258 5854 36260 5906
rect 36204 5852 36260 5854
rect 37884 10332 37940 10388
rect 39452 11394 39508 11396
rect 39452 11342 39454 11394
rect 39454 11342 39506 11394
rect 39506 11342 39508 11394
rect 39452 11340 39508 11342
rect 38556 10220 38612 10276
rect 38668 9772 38724 9828
rect 38556 9714 38612 9716
rect 38556 9662 38558 9714
rect 38558 9662 38610 9714
rect 38610 9662 38612 9714
rect 38556 9660 38612 9662
rect 40348 11452 40404 11508
rect 40460 11340 40516 11396
rect 39788 10668 39844 10724
rect 39676 10444 39732 10500
rect 39340 10220 39396 10276
rect 40460 9996 40516 10052
rect 40012 9826 40068 9828
rect 40012 9774 40014 9826
rect 40014 9774 40066 9826
rect 40066 9774 40068 9826
rect 40012 9772 40068 9774
rect 39788 9266 39844 9268
rect 39788 9214 39790 9266
rect 39790 9214 39842 9266
rect 39842 9214 39844 9266
rect 39788 9212 39844 9214
rect 41356 17612 41412 17668
rect 40796 16604 40852 16660
rect 40908 17388 40964 17444
rect 41132 17052 41188 17108
rect 41020 16882 41076 16884
rect 41020 16830 41022 16882
rect 41022 16830 41074 16882
rect 41074 16830 41076 16882
rect 41020 16828 41076 16830
rect 41692 17276 41748 17332
rect 41468 16604 41524 16660
rect 41356 16268 41412 16324
rect 41356 16098 41412 16100
rect 41356 16046 41358 16098
rect 41358 16046 41410 16098
rect 41410 16046 41412 16098
rect 41356 16044 41412 16046
rect 41468 15820 41524 15876
rect 41132 14924 41188 14980
rect 41132 14700 41188 14756
rect 41916 20188 41972 20244
rect 42476 21810 42532 21812
rect 42476 21758 42478 21810
rect 42478 21758 42530 21810
rect 42530 21758 42532 21810
rect 42476 21756 42532 21758
rect 43260 24834 43316 24836
rect 43260 24782 43262 24834
rect 43262 24782 43314 24834
rect 43314 24782 43316 24834
rect 43260 24780 43316 24782
rect 43148 24220 43204 24276
rect 42924 22988 42980 23044
rect 43036 24108 43092 24164
rect 43484 24498 43540 24500
rect 43484 24446 43486 24498
rect 43486 24446 43538 24498
rect 43538 24446 43540 24498
rect 43484 24444 43540 24446
rect 43036 21756 43092 21812
rect 42364 20914 42420 20916
rect 42364 20862 42366 20914
rect 42366 20862 42418 20914
rect 42418 20862 42420 20914
rect 42364 20860 42420 20862
rect 42700 20524 42756 20580
rect 42924 20018 42980 20020
rect 42924 19966 42926 20018
rect 42926 19966 42978 20018
rect 42978 19966 42980 20018
rect 42924 19964 42980 19966
rect 41916 17276 41972 17332
rect 41804 16882 41860 16884
rect 41804 16830 41806 16882
rect 41806 16830 41858 16882
rect 41858 16830 41860 16882
rect 41804 16828 41860 16830
rect 41916 16716 41972 16772
rect 41916 16322 41972 16324
rect 41916 16270 41918 16322
rect 41918 16270 41970 16322
rect 41970 16270 41972 16322
rect 41916 16268 41972 16270
rect 44268 23212 44324 23268
rect 43372 21698 43428 21700
rect 43372 21646 43374 21698
rect 43374 21646 43426 21698
rect 43426 21646 43428 21698
rect 43372 21644 43428 21646
rect 44604 23042 44660 23044
rect 44604 22990 44606 23042
rect 44606 22990 44658 23042
rect 44658 22990 44660 23042
rect 44604 22988 44660 22990
rect 43148 20860 43204 20916
rect 44044 20914 44100 20916
rect 44044 20862 44046 20914
rect 44046 20862 44098 20914
rect 44098 20862 44100 20914
rect 44044 20860 44100 20862
rect 44044 20412 44100 20468
rect 43708 20188 43764 20244
rect 43932 20188 43988 20244
rect 43260 18450 43316 18452
rect 43260 18398 43262 18450
rect 43262 18398 43314 18450
rect 43314 18398 43316 18450
rect 43260 18396 43316 18398
rect 42700 17666 42756 17668
rect 42700 17614 42702 17666
rect 42702 17614 42754 17666
rect 42754 17614 42756 17666
rect 42700 17612 42756 17614
rect 42588 16828 42644 16884
rect 42364 15874 42420 15876
rect 42364 15822 42366 15874
rect 42366 15822 42418 15874
rect 42418 15822 42420 15874
rect 42364 15820 42420 15822
rect 42364 15314 42420 15316
rect 42364 15262 42366 15314
rect 42366 15262 42418 15314
rect 42418 15262 42420 15314
rect 42364 15260 42420 15262
rect 43596 19852 43652 19908
rect 43708 19794 43764 19796
rect 43708 19742 43710 19794
rect 43710 19742 43762 19794
rect 43762 19742 43764 19794
rect 43708 19740 43764 19742
rect 43260 17500 43316 17556
rect 43372 17052 43428 17108
rect 43372 16882 43428 16884
rect 43372 16830 43374 16882
rect 43374 16830 43426 16882
rect 43426 16830 43428 16882
rect 43372 16828 43428 16830
rect 43036 15314 43092 15316
rect 43036 15262 43038 15314
rect 43038 15262 43090 15314
rect 43090 15262 43092 15314
rect 43036 15260 43092 15262
rect 41468 14028 41524 14084
rect 41804 14306 41860 14308
rect 41804 14254 41806 14306
rect 41806 14254 41858 14306
rect 41858 14254 41860 14306
rect 41804 14252 41860 14254
rect 41692 12066 41748 12068
rect 41692 12014 41694 12066
rect 41694 12014 41746 12066
rect 41746 12014 41748 12066
rect 41692 12012 41748 12014
rect 41132 11506 41188 11508
rect 41132 11454 41134 11506
rect 41134 11454 41186 11506
rect 41186 11454 41188 11506
rect 41132 11452 41188 11454
rect 41916 13356 41972 13412
rect 42140 14812 42196 14868
rect 44044 18562 44100 18564
rect 44044 18510 44046 18562
rect 44046 18510 44098 18562
rect 44098 18510 44100 18562
rect 44044 18508 44100 18510
rect 43820 16994 43876 16996
rect 43820 16942 43822 16994
rect 43822 16942 43874 16994
rect 43874 16942 43876 16994
rect 43820 16940 43876 16942
rect 43484 14812 43540 14868
rect 42364 14700 42420 14756
rect 42812 14418 42868 14420
rect 42812 14366 42814 14418
rect 42814 14366 42866 14418
rect 42866 14366 42868 14418
rect 42812 14364 42868 14366
rect 42252 14028 42308 14084
rect 43148 14588 43204 14644
rect 43148 14252 43204 14308
rect 43484 13858 43540 13860
rect 43484 13806 43486 13858
rect 43486 13806 43538 13858
rect 43538 13806 43540 13858
rect 43484 13804 43540 13806
rect 43820 14642 43876 14644
rect 43820 14590 43822 14642
rect 43822 14590 43874 14642
rect 43874 14590 43876 14642
rect 43820 14588 43876 14590
rect 44268 17388 44324 17444
rect 42028 12962 42084 12964
rect 42028 12910 42030 12962
rect 42030 12910 42082 12962
rect 42082 12910 42084 12962
rect 42028 12908 42084 12910
rect 41804 11394 41860 11396
rect 41804 11342 41806 11394
rect 41806 11342 41858 11394
rect 41858 11342 41860 11394
rect 41804 11340 41860 11342
rect 40684 9660 40740 9716
rect 40460 9266 40516 9268
rect 40460 9214 40462 9266
rect 40462 9214 40514 9266
rect 40514 9214 40516 9266
rect 40460 9212 40516 9214
rect 37436 6524 37492 6580
rect 37324 6466 37380 6468
rect 37324 6414 37326 6466
rect 37326 6414 37378 6466
rect 37378 6414 37380 6466
rect 37324 6412 37380 6414
rect 36876 5852 36932 5908
rect 37660 5794 37716 5796
rect 37660 5742 37662 5794
rect 37662 5742 37714 5794
rect 37714 5742 37716 5794
rect 37660 5740 37716 5742
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35644 5010 35700 5012
rect 35644 4958 35646 5010
rect 35646 4958 35698 5010
rect 35698 4958 35700 5010
rect 35644 4956 35700 4958
rect 35084 4508 35140 4564
rect 39116 7980 39172 8036
rect 39004 7420 39060 7476
rect 38108 6690 38164 6692
rect 38108 6638 38110 6690
rect 38110 6638 38162 6690
rect 38162 6638 38164 6690
rect 38108 6636 38164 6638
rect 38668 6690 38724 6692
rect 38668 6638 38670 6690
rect 38670 6638 38722 6690
rect 38722 6638 38724 6690
rect 38668 6636 38724 6638
rect 38444 6466 38500 6468
rect 38444 6414 38446 6466
rect 38446 6414 38498 6466
rect 38498 6414 38500 6466
rect 38444 6412 38500 6414
rect 38444 5906 38500 5908
rect 38444 5854 38446 5906
rect 38446 5854 38498 5906
rect 38498 5854 38500 5906
rect 38444 5852 38500 5854
rect 37884 4732 37940 4788
rect 35532 4508 35588 4564
rect 38668 5122 38724 5124
rect 38668 5070 38670 5122
rect 38670 5070 38722 5122
rect 38722 5070 38724 5122
rect 38668 5068 38724 5070
rect 39676 5906 39732 5908
rect 39676 5854 39678 5906
rect 39678 5854 39730 5906
rect 39730 5854 39732 5906
rect 39676 5852 39732 5854
rect 40012 5852 40068 5908
rect 39452 5740 39508 5796
rect 39788 5516 39844 5572
rect 39452 5292 39508 5348
rect 39004 5068 39060 5124
rect 39116 5180 39172 5236
rect 38444 4508 38500 4564
rect 35308 4396 35364 4452
rect 34972 4284 35028 4340
rect 34412 4226 34468 4228
rect 34412 4174 34414 4226
rect 34414 4174 34466 4226
rect 34466 4174 34468 4226
rect 34412 4172 34468 4174
rect 39004 4450 39060 4452
rect 39004 4398 39006 4450
rect 39006 4398 39058 4450
rect 39058 4398 39060 4450
rect 39004 4396 39060 4398
rect 38108 4226 38164 4228
rect 38108 4174 38110 4226
rect 38110 4174 38162 4226
rect 38162 4174 38164 4226
rect 38108 4172 38164 4174
rect 35868 4114 35924 4116
rect 35868 4062 35870 4114
rect 35870 4062 35922 4114
rect 35922 4062 35924 4114
rect 35868 4060 35924 4062
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 39340 5068 39396 5124
rect 40348 5852 40404 5908
rect 39564 4562 39620 4564
rect 39564 4510 39566 4562
rect 39566 4510 39618 4562
rect 39618 4510 39620 4562
rect 39564 4508 39620 4510
rect 40012 5404 40068 5460
rect 40572 5516 40628 5572
rect 40796 5346 40852 5348
rect 40796 5294 40798 5346
rect 40798 5294 40850 5346
rect 40850 5294 40852 5346
rect 40796 5292 40852 5294
rect 40460 5068 40516 5124
rect 40460 4620 40516 4676
rect 41468 10780 41524 10836
rect 41692 11170 41748 11172
rect 41692 11118 41694 11170
rect 41694 11118 41746 11170
rect 41746 11118 41748 11170
rect 41692 11116 41748 11118
rect 41356 9714 41412 9716
rect 41356 9662 41358 9714
rect 41358 9662 41410 9714
rect 41410 9662 41412 9714
rect 41356 9660 41412 9662
rect 42028 11340 42084 11396
rect 42252 11228 42308 11284
rect 42140 10892 42196 10948
rect 42364 10610 42420 10612
rect 42364 10558 42366 10610
rect 42366 10558 42418 10610
rect 42418 10558 42420 10610
rect 42364 10556 42420 10558
rect 43036 13356 43092 13412
rect 43484 13580 43540 13636
rect 42588 12962 42644 12964
rect 42588 12910 42590 12962
rect 42590 12910 42642 12962
rect 42642 12910 42644 12962
rect 42588 12908 42644 12910
rect 42588 12066 42644 12068
rect 42588 12014 42590 12066
rect 42590 12014 42642 12066
rect 42642 12014 42644 12066
rect 42588 12012 42644 12014
rect 42924 12124 42980 12180
rect 43372 12178 43428 12180
rect 43372 12126 43374 12178
rect 43374 12126 43426 12178
rect 43426 12126 43428 12178
rect 43372 12124 43428 12126
rect 44044 12066 44100 12068
rect 44044 12014 44046 12066
rect 44046 12014 44098 12066
rect 44098 12014 44100 12066
rect 44044 12012 44100 12014
rect 43372 11394 43428 11396
rect 43372 11342 43374 11394
rect 43374 11342 43426 11394
rect 43426 11342 43428 11394
rect 43372 11340 43428 11342
rect 43708 11394 43764 11396
rect 43708 11342 43710 11394
rect 43710 11342 43762 11394
rect 43762 11342 43764 11394
rect 43708 11340 43764 11342
rect 43932 11282 43988 11284
rect 43932 11230 43934 11282
rect 43934 11230 43986 11282
rect 43986 11230 43988 11282
rect 43932 11228 43988 11230
rect 42924 11116 42980 11172
rect 43036 10610 43092 10612
rect 43036 10558 43038 10610
rect 43038 10558 43090 10610
rect 43090 10558 43092 10610
rect 43036 10556 43092 10558
rect 41244 7308 41300 7364
rect 41468 8258 41524 8260
rect 41468 8206 41470 8258
rect 41470 8206 41522 8258
rect 41522 8206 41524 8258
rect 41468 8204 41524 8206
rect 43820 9772 43876 9828
rect 42588 9660 42644 9716
rect 42476 8258 42532 8260
rect 42476 8206 42478 8258
rect 42478 8206 42530 8258
rect 42530 8206 42532 8258
rect 42476 8204 42532 8206
rect 42812 8316 42868 8372
rect 43820 8988 43876 9044
rect 43148 8370 43204 8372
rect 43148 8318 43150 8370
rect 43150 8318 43202 8370
rect 43202 8318 43204 8370
rect 43148 8316 43204 8318
rect 44716 18508 44772 18564
rect 44604 16940 44660 16996
rect 47068 25452 47124 25508
rect 55580 25506 55636 25508
rect 55580 25454 55582 25506
rect 55582 25454 55634 25506
rect 55634 25454 55636 25506
rect 55580 25452 55636 25454
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 58268 26236 58324 26292
rect 58156 25564 58212 25620
rect 57932 24892 57988 24948
rect 46172 24444 46228 24500
rect 45500 23714 45556 23716
rect 45500 23662 45502 23714
rect 45502 23662 45554 23714
rect 45554 23662 45556 23714
rect 45500 23660 45556 23662
rect 44940 23266 44996 23268
rect 44940 23214 44942 23266
rect 44942 23214 44994 23266
rect 44994 23214 44996 23266
rect 44940 23212 44996 23214
rect 45388 22988 45444 23044
rect 44940 22370 44996 22372
rect 44940 22318 44942 22370
rect 44942 22318 44994 22370
rect 44994 22318 44996 22370
rect 44940 22316 44996 22318
rect 45948 23548 46004 23604
rect 50092 23884 50148 23940
rect 55580 23938 55636 23940
rect 55580 23886 55582 23938
rect 55582 23886 55634 23938
rect 55634 23886 55636 23938
rect 55580 23884 55636 23886
rect 47292 23548 47348 23604
rect 46172 23212 46228 23268
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 57932 23548 57988 23604
rect 50764 23492 50820 23494
rect 47852 23100 47908 23156
rect 48748 23100 48804 23156
rect 45276 22428 45332 22484
rect 45052 22204 45108 22260
rect 46844 23042 46900 23044
rect 46844 22990 46846 23042
rect 46846 22990 46898 23042
rect 46898 22990 46900 23042
rect 46844 22988 46900 22990
rect 45724 22370 45780 22372
rect 45724 22318 45726 22370
rect 45726 22318 45778 22370
rect 45778 22318 45780 22370
rect 45724 22316 45780 22318
rect 49084 23154 49140 23156
rect 49084 23102 49086 23154
rect 49086 23102 49138 23154
rect 49138 23102 49140 23154
rect 49084 23100 49140 23102
rect 48860 23042 48916 23044
rect 48860 22990 48862 23042
rect 48862 22990 48914 23042
rect 48914 22990 48916 23042
rect 48860 22988 48916 22990
rect 51100 22316 51156 22372
rect 46172 22258 46228 22260
rect 46172 22206 46174 22258
rect 46174 22206 46226 22258
rect 46226 22206 46228 22258
rect 46172 22204 46228 22206
rect 44940 20188 44996 20244
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 55580 22370 55636 22372
rect 55580 22318 55582 22370
rect 55582 22318 55634 22370
rect 55634 22318 55636 22370
rect 55580 22316 55636 22318
rect 46172 20690 46228 20692
rect 46172 20638 46174 20690
rect 46174 20638 46226 20690
rect 46226 20638 46228 20690
rect 46172 20636 46228 20638
rect 47292 20860 47348 20916
rect 46956 20748 47012 20804
rect 45612 20412 45668 20468
rect 45948 20076 46004 20132
rect 45948 19906 46004 19908
rect 45948 19854 45950 19906
rect 45950 19854 46002 19906
rect 46002 19854 46004 19906
rect 45948 19852 46004 19854
rect 45388 16268 45444 16324
rect 45724 16156 45780 16212
rect 46284 19740 46340 19796
rect 48636 20914 48692 20916
rect 48636 20862 48638 20914
rect 48638 20862 48690 20914
rect 48690 20862 48692 20914
rect 48636 20860 48692 20862
rect 49532 20914 49588 20916
rect 49532 20862 49534 20914
rect 49534 20862 49586 20914
rect 49586 20862 49588 20914
rect 49532 20860 49588 20862
rect 47964 20802 48020 20804
rect 47964 20750 47966 20802
rect 47966 20750 48018 20802
rect 48018 20750 48020 20802
rect 47964 20748 48020 20750
rect 58156 22204 58212 22260
rect 57932 21532 57988 21588
rect 48860 20636 48916 20692
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 58156 20242 58212 20244
rect 58156 20190 58158 20242
rect 58158 20190 58210 20242
rect 58210 20190 58212 20242
rect 58156 20188 58212 20190
rect 47068 20076 47124 20132
rect 49196 20130 49252 20132
rect 49196 20078 49198 20130
rect 49198 20078 49250 20130
rect 49250 20078 49252 20130
rect 49196 20076 49252 20078
rect 47964 19740 48020 19796
rect 48972 19740 49028 19796
rect 49308 19740 49364 19796
rect 49532 19122 49588 19124
rect 49532 19070 49534 19122
rect 49534 19070 49586 19122
rect 49586 19070 49588 19122
rect 49532 19068 49588 19070
rect 46060 18396 46116 18452
rect 45948 18284 46004 18340
rect 48748 18396 48804 18452
rect 45948 15260 46004 15316
rect 45612 15036 45668 15092
rect 45052 14418 45108 14420
rect 45052 14366 45054 14418
rect 45054 14366 45106 14418
rect 45106 14366 45108 14418
rect 45052 14364 45108 14366
rect 44940 14306 44996 14308
rect 44940 14254 44942 14306
rect 44942 14254 44994 14306
rect 44994 14254 44996 14306
rect 44940 14252 44996 14254
rect 45164 13970 45220 13972
rect 45164 13918 45166 13970
rect 45166 13918 45218 13970
rect 45218 13918 45220 13970
rect 45164 13916 45220 13918
rect 44828 13858 44884 13860
rect 44828 13806 44830 13858
rect 44830 13806 44882 13858
rect 44882 13806 44884 13858
rect 44828 13804 44884 13806
rect 45500 13858 45556 13860
rect 45500 13806 45502 13858
rect 45502 13806 45554 13858
rect 45554 13806 45556 13858
rect 45500 13804 45556 13806
rect 45388 13634 45444 13636
rect 45388 13582 45390 13634
rect 45390 13582 45442 13634
rect 45442 13582 45444 13634
rect 45388 13580 45444 13582
rect 45836 14812 45892 14868
rect 46172 14588 46228 14644
rect 45724 14306 45780 14308
rect 45724 14254 45726 14306
rect 45726 14254 45778 14306
rect 45778 14254 45780 14306
rect 45724 14252 45780 14254
rect 45836 13746 45892 13748
rect 45836 13694 45838 13746
rect 45838 13694 45890 13746
rect 45890 13694 45892 13746
rect 45836 13692 45892 13694
rect 46172 14306 46228 14308
rect 46172 14254 46174 14306
rect 46174 14254 46226 14306
rect 46226 14254 46228 14306
rect 46172 14252 46228 14254
rect 46172 13580 46228 13636
rect 45612 13468 45668 13524
rect 46508 17666 46564 17668
rect 46508 17614 46510 17666
rect 46510 17614 46562 17666
rect 46562 17614 46564 17666
rect 46508 17612 46564 17614
rect 47068 17666 47124 17668
rect 47068 17614 47070 17666
rect 47070 17614 47122 17666
rect 47122 17614 47124 17666
rect 47068 17612 47124 17614
rect 47292 17612 47348 17668
rect 46844 16940 46900 16996
rect 46956 17500 47012 17556
rect 47516 17724 47572 17780
rect 47404 17500 47460 17556
rect 49644 18450 49700 18452
rect 49644 18398 49646 18450
rect 49646 18398 49698 18450
rect 49698 18398 49700 18450
rect 49644 18396 49700 18398
rect 49532 17724 49588 17780
rect 48076 17666 48132 17668
rect 48076 17614 48078 17666
rect 48078 17614 48130 17666
rect 48130 17614 48132 17666
rect 48076 17612 48132 17614
rect 48636 17666 48692 17668
rect 48636 17614 48638 17666
rect 48638 17614 48690 17666
rect 48690 17614 48692 17666
rect 48636 17612 48692 17614
rect 49196 17666 49252 17668
rect 49196 17614 49198 17666
rect 49198 17614 49250 17666
rect 49250 17614 49252 17666
rect 49196 17612 49252 17614
rect 50428 19180 50484 19236
rect 50092 17500 50148 17556
rect 50204 19122 50260 19124
rect 50204 19070 50206 19122
rect 50206 19070 50258 19122
rect 50258 19070 50260 19122
rect 50204 19068 50260 19070
rect 51436 19234 51492 19236
rect 51436 19182 51438 19234
rect 51438 19182 51490 19234
rect 51490 19182 51492 19234
rect 51436 19180 51492 19182
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 50316 18338 50372 18340
rect 50316 18286 50318 18338
rect 50318 18286 50370 18338
rect 50370 18286 50372 18338
rect 50316 18284 50372 18286
rect 51660 18284 51716 18340
rect 50204 17612 50260 17668
rect 51324 17666 51380 17668
rect 51324 17614 51326 17666
rect 51326 17614 51378 17666
rect 51378 17614 51380 17666
rect 51324 17612 51380 17614
rect 50652 17554 50708 17556
rect 50652 17502 50654 17554
rect 50654 17502 50706 17554
rect 50706 17502 50708 17554
rect 50652 17500 50708 17502
rect 51100 17554 51156 17556
rect 51100 17502 51102 17554
rect 51102 17502 51154 17554
rect 51154 17502 51156 17554
rect 51100 17500 51156 17502
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 47516 16828 47572 16884
rect 58156 18844 58212 18900
rect 57932 18172 57988 18228
rect 53004 17612 53060 17668
rect 55580 17666 55636 17668
rect 55580 17614 55582 17666
rect 55582 17614 55634 17666
rect 55634 17614 55636 17666
rect 55580 17612 55636 17614
rect 46844 16658 46900 16660
rect 46844 16606 46846 16658
rect 46846 16606 46898 16658
rect 46898 16606 46900 16658
rect 46844 16604 46900 16606
rect 47628 16604 47684 16660
rect 46396 14588 46452 14644
rect 46508 13916 46564 13972
rect 46620 14812 46676 14868
rect 46396 13746 46452 13748
rect 46396 13694 46398 13746
rect 46398 13694 46450 13746
rect 46450 13694 46452 13746
rect 46396 13692 46452 13694
rect 44492 12178 44548 12180
rect 44492 12126 44494 12178
rect 44494 12126 44546 12178
rect 44546 12126 44548 12178
rect 44492 12124 44548 12126
rect 44156 9826 44212 9828
rect 44156 9774 44158 9826
rect 44158 9774 44210 9826
rect 44210 9774 44212 9826
rect 44156 9772 44212 9774
rect 45388 9996 45444 10052
rect 50204 16156 50260 16212
rect 50092 16044 50148 16100
rect 49868 15874 49924 15876
rect 49868 15822 49870 15874
rect 49870 15822 49922 15874
rect 49922 15822 49924 15874
rect 49868 15820 49924 15822
rect 47068 15314 47124 15316
rect 47068 15262 47070 15314
rect 47070 15262 47122 15314
rect 47122 15262 47124 15314
rect 47068 15260 47124 15262
rect 48300 15426 48356 15428
rect 48300 15374 48302 15426
rect 48302 15374 48354 15426
rect 48354 15374 48356 15426
rect 48300 15372 48356 15374
rect 47068 14252 47124 14308
rect 47404 13970 47460 13972
rect 47404 13918 47406 13970
rect 47406 13918 47458 13970
rect 47458 13918 47460 13970
rect 47404 13916 47460 13918
rect 46732 13858 46788 13860
rect 46732 13806 46734 13858
rect 46734 13806 46786 13858
rect 46786 13806 46788 13858
rect 46732 13804 46788 13806
rect 47292 13746 47348 13748
rect 47292 13694 47294 13746
rect 47294 13694 47346 13746
rect 47346 13694 47348 13746
rect 47292 13692 47348 13694
rect 49532 13692 49588 13748
rect 46844 13020 46900 13076
rect 47292 13468 47348 13524
rect 46620 12012 46676 12068
rect 46956 11340 47012 11396
rect 51884 16828 51940 16884
rect 53116 16882 53172 16884
rect 53116 16830 53118 16882
rect 53118 16830 53170 16882
rect 53170 16830 53172 16882
rect 53116 16828 53172 16830
rect 51212 16210 51268 16212
rect 51212 16158 51214 16210
rect 51214 16158 51266 16210
rect 51266 16158 51268 16210
rect 51212 16156 51268 16158
rect 57932 16716 57988 16772
rect 50876 16098 50932 16100
rect 50876 16046 50878 16098
rect 50878 16046 50930 16098
rect 50930 16046 50932 16098
rect 50876 16044 50932 16046
rect 51548 15986 51604 15988
rect 51548 15934 51550 15986
rect 51550 15934 51602 15986
rect 51602 15934 51604 15986
rect 51548 15932 51604 15934
rect 50988 15820 51044 15876
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 51100 15426 51156 15428
rect 51100 15374 51102 15426
rect 51102 15374 51154 15426
rect 51154 15374 51156 15426
rect 51100 15372 51156 15374
rect 51324 15148 51380 15204
rect 58156 16156 58212 16212
rect 53004 16044 53060 16100
rect 52668 15986 52724 15988
rect 52668 15934 52670 15986
rect 52670 15934 52722 15986
rect 52722 15934 52724 15986
rect 52668 15932 52724 15934
rect 55580 16098 55636 16100
rect 55580 16046 55582 16098
rect 55582 16046 55634 16098
rect 55634 16046 55636 16098
rect 55580 16044 55636 16046
rect 57932 15484 57988 15540
rect 52332 15372 52388 15428
rect 51884 15202 51940 15204
rect 51884 15150 51886 15202
rect 51886 15150 51938 15202
rect 51938 15150 51940 15202
rect 51884 15148 51940 15150
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 48972 13074 49028 13076
rect 48972 13022 48974 13074
rect 48974 13022 49026 13074
rect 49026 13022 49028 13074
rect 48972 13020 49028 13022
rect 50092 13020 50148 13076
rect 49196 12962 49252 12964
rect 49196 12910 49198 12962
rect 49198 12910 49250 12962
rect 49250 12910 49252 12962
rect 49196 12908 49252 12910
rect 47516 12290 47572 12292
rect 47516 12238 47518 12290
rect 47518 12238 47570 12290
rect 47570 12238 47572 12290
rect 47516 12236 47572 12238
rect 49196 12236 49252 12292
rect 50204 12908 50260 12964
rect 53340 14476 53396 14532
rect 55580 14530 55636 14532
rect 55580 14478 55582 14530
rect 55582 14478 55634 14530
rect 55634 14478 55636 14530
rect 55580 14476 55636 14478
rect 52220 13746 52276 13748
rect 52220 13694 52222 13746
rect 52222 13694 52274 13746
rect 52274 13694 52276 13746
rect 52220 13692 52276 13694
rect 58156 13468 58212 13524
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 58156 12124 58212 12180
rect 47516 11394 47572 11396
rect 47516 11342 47518 11394
rect 47518 11342 47570 11394
rect 47570 11342 47572 11394
rect 47516 11340 47572 11342
rect 47852 11170 47908 11172
rect 47852 11118 47854 11170
rect 47854 11118 47906 11170
rect 47906 11118 47908 11170
rect 47852 11116 47908 11118
rect 45052 9826 45108 9828
rect 45052 9774 45054 9826
rect 45054 9774 45106 9826
rect 45106 9774 45108 9826
rect 45052 9772 45108 9774
rect 45388 9772 45444 9828
rect 48972 11116 49028 11172
rect 46732 10610 46788 10612
rect 46732 10558 46734 10610
rect 46734 10558 46786 10610
rect 46786 10558 46788 10610
rect 46732 10556 46788 10558
rect 47180 10556 47236 10612
rect 46284 9938 46340 9940
rect 46284 9886 46286 9938
rect 46286 9886 46338 9938
rect 46338 9886 46340 9938
rect 46284 9884 46340 9886
rect 47068 9938 47124 9940
rect 47068 9886 47070 9938
rect 47070 9886 47122 9938
rect 47122 9886 47124 9938
rect 47068 9884 47124 9886
rect 46508 9826 46564 9828
rect 46508 9774 46510 9826
rect 46510 9774 46562 9826
rect 46562 9774 46564 9826
rect 46508 9772 46564 9774
rect 47628 10610 47684 10612
rect 47628 10558 47630 10610
rect 47630 10558 47682 10610
rect 47682 10558 47684 10610
rect 47628 10556 47684 10558
rect 48860 10610 48916 10612
rect 48860 10558 48862 10610
rect 48862 10558 48914 10610
rect 48914 10558 48916 10610
rect 48860 10556 48916 10558
rect 49084 9602 49140 9604
rect 49084 9550 49086 9602
rect 49086 9550 49138 9602
rect 49138 9550 49140 9602
rect 49084 9548 49140 9550
rect 49980 9548 50036 9604
rect 47852 9100 47908 9156
rect 44940 9042 44996 9044
rect 44940 8990 44942 9042
rect 44942 8990 44994 9042
rect 44994 8990 44996 9042
rect 44940 8988 44996 8990
rect 44268 8764 44324 8820
rect 44716 8818 44772 8820
rect 44716 8766 44718 8818
rect 44718 8766 44770 8818
rect 44770 8766 44772 8818
rect 44716 8764 44772 8766
rect 43932 8316 43988 8372
rect 43036 8204 43092 8260
rect 42700 7756 42756 7812
rect 43372 7980 43428 8036
rect 42028 7644 42084 7700
rect 42252 7474 42308 7476
rect 42252 7422 42254 7474
rect 42254 7422 42306 7474
rect 42306 7422 42308 7474
rect 42252 7420 42308 7422
rect 41468 6300 41524 6356
rect 41244 5906 41300 5908
rect 41244 5854 41246 5906
rect 41246 5854 41298 5906
rect 41298 5854 41300 5906
rect 41244 5852 41300 5854
rect 41468 5516 41524 5572
rect 45388 8316 45444 8372
rect 45164 8258 45220 8260
rect 45164 8206 45166 8258
rect 45166 8206 45218 8258
rect 45218 8206 45220 8258
rect 45164 8204 45220 8206
rect 45500 8204 45556 8260
rect 45500 7868 45556 7924
rect 42812 6076 42868 6132
rect 42140 5628 42196 5684
rect 41916 5516 41972 5572
rect 42924 5682 42980 5684
rect 42924 5630 42926 5682
rect 42926 5630 42978 5682
rect 42978 5630 42980 5682
rect 42924 5628 42980 5630
rect 42364 5404 42420 5460
rect 43148 5906 43204 5908
rect 43148 5854 43150 5906
rect 43150 5854 43202 5906
rect 43202 5854 43204 5906
rect 43148 5852 43204 5854
rect 42140 5180 42196 5236
rect 42140 5010 42196 5012
rect 42140 4958 42142 5010
rect 42142 4958 42194 5010
rect 42194 4958 42196 5010
rect 42140 4956 42196 4958
rect 41916 4844 41972 4900
rect 44268 6130 44324 6132
rect 44268 6078 44270 6130
rect 44270 6078 44322 6130
rect 44322 6078 44324 6130
rect 44268 6076 44324 6078
rect 43708 5682 43764 5684
rect 43708 5630 43710 5682
rect 43710 5630 43762 5682
rect 43762 5630 43764 5682
rect 43708 5628 43764 5630
rect 43036 4956 43092 5012
rect 42812 4450 42868 4452
rect 42812 4398 42814 4450
rect 42814 4398 42866 4450
rect 42866 4398 42868 4450
rect 42812 4396 42868 4398
rect 44604 5906 44660 5908
rect 44604 5854 44606 5906
rect 44606 5854 44658 5906
rect 44658 5854 44660 5906
rect 44604 5852 44660 5854
rect 46172 7868 46228 7924
rect 47068 7362 47124 7364
rect 47068 7310 47070 7362
rect 47070 7310 47122 7362
rect 47122 7310 47124 7362
rect 47068 7308 47124 7310
rect 49084 9154 49140 9156
rect 49084 9102 49086 9154
rect 49086 9102 49138 9154
rect 49138 9102 49140 9154
rect 49084 9100 49140 9102
rect 48188 8876 48244 8932
rect 49196 8930 49252 8932
rect 49196 8878 49198 8930
rect 49198 8878 49250 8930
rect 49250 8878 49252 8930
rect 49196 8876 49252 8878
rect 48300 7308 48356 7364
rect 49084 7420 49140 7476
rect 49532 8988 49588 9044
rect 57932 11506 57988 11508
rect 57932 11454 57934 11506
rect 57934 11454 57986 11506
rect 57986 11454 57988 11506
rect 57932 11452 57988 11454
rect 51660 11340 51716 11396
rect 55580 11394 55636 11396
rect 55580 11342 55582 11394
rect 55582 11342 55634 11394
rect 55634 11342 55636 11394
rect 55580 11340 55636 11342
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 58156 10780 58212 10836
rect 57708 10108 57764 10164
rect 51436 9548 51492 9604
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 58156 9436 58212 9492
rect 50204 8988 50260 9044
rect 50652 8988 50708 9044
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 50876 7474 50932 7476
rect 50876 7422 50878 7474
rect 50878 7422 50930 7474
rect 50930 7422 50932 7474
rect 50876 7420 50932 7422
rect 57932 8370 57988 8372
rect 57932 8318 57934 8370
rect 57934 8318 57986 8370
rect 57986 8318 57988 8370
rect 57932 8316 57988 8318
rect 51996 8204 52052 8260
rect 55580 8258 55636 8260
rect 55580 8206 55582 8258
rect 55582 8206 55634 8258
rect 55634 8206 55636 8258
rect 55580 8204 55636 8206
rect 58156 8092 58212 8148
rect 49420 7362 49476 7364
rect 49420 7310 49422 7362
rect 49422 7310 49474 7362
rect 49474 7310 49476 7362
rect 49420 7308 49476 7310
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 48748 6018 48804 6020
rect 48748 5966 48750 6018
rect 48750 5966 48802 6018
rect 48802 5966 48804 6018
rect 48748 5964 48804 5966
rect 46060 5852 46116 5908
rect 46732 5906 46788 5908
rect 46732 5854 46734 5906
rect 46734 5854 46786 5906
rect 46786 5854 46788 5906
rect 46732 5852 46788 5854
rect 47628 5906 47684 5908
rect 47628 5854 47630 5906
rect 47630 5854 47682 5906
rect 47682 5854 47684 5906
rect 47628 5852 47684 5854
rect 48412 5852 48468 5908
rect 44380 5682 44436 5684
rect 44380 5630 44382 5682
rect 44382 5630 44434 5682
rect 44434 5630 44436 5682
rect 44380 5628 44436 5630
rect 44380 5180 44436 5236
rect 45164 5068 45220 5124
rect 44044 5010 44100 5012
rect 44044 4958 44046 5010
rect 44046 4958 44098 5010
rect 44098 4958 44100 5010
rect 44044 4956 44100 4958
rect 44156 4898 44212 4900
rect 44156 4846 44158 4898
rect 44158 4846 44210 4898
rect 44210 4846 44212 4898
rect 44156 4844 44212 4846
rect 43708 4060 43764 4116
rect 41132 3276 41188 3332
rect 42364 3612 42420 3668
rect 30492 1596 30548 1652
rect 46396 5516 46452 5572
rect 46508 5740 46564 5796
rect 46060 5122 46116 5124
rect 46060 5070 46062 5122
rect 46062 5070 46114 5122
rect 46114 5070 46116 5122
rect 46060 5068 46116 5070
rect 47292 5794 47348 5796
rect 47292 5742 47294 5794
rect 47294 5742 47346 5794
rect 47346 5742 47348 5794
rect 47292 5740 47348 5742
rect 48188 5682 48244 5684
rect 48188 5630 48190 5682
rect 48190 5630 48242 5682
rect 48242 5630 48244 5682
rect 48188 5628 48244 5630
rect 47852 5516 47908 5572
rect 46732 5234 46788 5236
rect 46732 5182 46734 5234
rect 46734 5182 46786 5234
rect 46786 5182 46788 5234
rect 46732 5180 46788 5182
rect 48076 5234 48132 5236
rect 48076 5182 48078 5234
rect 48078 5182 48130 5234
rect 48130 5182 48132 5234
rect 48076 5180 48132 5182
rect 47068 5122 47124 5124
rect 47068 5070 47070 5122
rect 47070 5070 47122 5122
rect 47122 5070 47124 5122
rect 47068 5068 47124 5070
rect 45388 4844 45444 4900
rect 45276 4620 45332 4676
rect 48860 5852 48916 5908
rect 49420 5964 49476 6020
rect 49644 5906 49700 5908
rect 49644 5854 49646 5906
rect 49646 5854 49698 5906
rect 49698 5854 49700 5906
rect 49644 5852 49700 5854
rect 50092 5628 50148 5684
rect 50092 5122 50148 5124
rect 50092 5070 50094 5122
rect 50094 5070 50146 5122
rect 50146 5070 50148 5122
rect 50092 5068 50148 5070
rect 48972 4956 49028 5012
rect 47404 4620 47460 4676
rect 44940 4114 44996 4116
rect 44940 4062 44942 4114
rect 44942 4062 44994 4114
rect 44994 4062 44996 4114
rect 44940 4060 44996 4062
rect 47180 3948 47236 4004
rect 44604 3666 44660 3668
rect 44604 3614 44606 3666
rect 44606 3614 44658 3666
rect 44658 3614 44660 3666
rect 44604 3612 44660 3614
rect 49084 4620 49140 4676
rect 49644 4620 49700 4676
rect 50764 4898 50820 4900
rect 50764 4846 50766 4898
rect 50766 4846 50818 4898
rect 50818 4846 50820 4898
rect 50764 4844 50820 4846
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 51212 5068 51268 5124
rect 51324 5010 51380 5012
rect 51324 4958 51326 5010
rect 51326 4958 51378 5010
rect 51378 4958 51380 5010
rect 51324 4956 51380 4958
rect 51436 4844 51492 4900
rect 48860 3948 48916 4004
rect 51100 4060 51156 4116
rect 50428 3612 50484 3668
rect 46396 3388 46452 3444
rect 48972 3442 49028 3444
rect 48972 3390 48974 3442
rect 48974 3390 49026 3442
rect 49026 3390 49028 3442
rect 48972 3388 49028 3390
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
rect 52332 4114 52388 4116
rect 52332 4062 52334 4114
rect 52334 4062 52386 4114
rect 52386 4062 52388 4114
rect 52332 4060 52388 4062
rect 52220 3666 52276 3668
rect 52220 3614 52222 3666
rect 52222 3614 52274 3666
rect 52274 3614 52276 3666
rect 52220 3612 52276 3614
rect 52444 3276 52500 3332
rect 54124 3330 54180 3332
rect 54124 3278 54126 3330
rect 54126 3278 54178 3330
rect 54178 3278 54180 3330
rect 54124 3276 54180 3278
<< metal3 >>
rect 20514 57820 20524 57876
rect 20580 57820 26684 57876
rect 26740 57820 26750 57876
rect 15026 57708 15036 57764
rect 15092 57708 36316 57764
rect 36372 57708 36382 57764
rect 12002 57596 12012 57652
rect 12068 57596 30604 57652
rect 30660 57596 30670 57652
rect 24994 57484 25004 57540
rect 25060 57484 38556 57540
rect 38612 57484 38622 57540
rect 22978 57372 22988 57428
rect 23044 57372 40572 57428
rect 40628 57372 40638 57428
rect 21074 57260 21084 57316
rect 21140 57260 27580 57316
rect 27636 57260 27646 57316
rect 16370 57148 16380 57204
rect 16436 57148 26460 57204
rect 26516 57148 26526 57204
rect 26674 57148 26684 57204
rect 26740 57148 40460 57204
rect 40516 57148 40526 57204
rect 21410 56700 21420 56756
rect 21476 56700 37100 56756
rect 37156 56700 37166 56756
rect 18274 56588 18284 56644
rect 18340 56588 19628 56644
rect 19684 56588 27020 56644
rect 27076 56588 27086 56644
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 20188 56364 24780 56420
rect 24836 56364 24846 56420
rect 20188 56308 20244 56364
rect 18162 56252 18172 56308
rect 18228 56252 20244 56308
rect 23314 56252 23324 56308
rect 23380 56252 34300 56308
rect 34356 56252 34366 56308
rect 45714 56252 45724 56308
rect 45780 56252 48412 56308
rect 48468 56252 48478 56308
rect 13794 56140 13804 56196
rect 13860 56140 15596 56196
rect 15652 56140 15662 56196
rect 17826 56140 17836 56196
rect 17892 56140 19180 56196
rect 19236 56140 19246 56196
rect 20962 56140 20972 56196
rect 21028 56140 21868 56196
rect 21924 56140 21934 56196
rect 22642 56140 22652 56196
rect 22708 56140 24668 56196
rect 24724 56140 25564 56196
rect 25620 56140 25630 56196
rect 28690 56140 28700 56196
rect 28756 56140 37436 56196
rect 37492 56140 37502 56196
rect 12562 56028 12572 56084
rect 12628 56028 20188 56084
rect 20244 56028 20254 56084
rect 20402 56028 20412 56084
rect 20468 56028 21308 56084
rect 21364 56028 21374 56084
rect 23538 56028 23548 56084
rect 23604 56028 30716 56084
rect 30772 56028 36988 56084
rect 37044 56028 37054 56084
rect 41682 56028 41692 56084
rect 41748 56028 42588 56084
rect 42644 56028 42654 56084
rect 46498 56028 46508 56084
rect 46564 56028 47404 56084
rect 47460 56028 47470 56084
rect 52994 56028 53004 56084
rect 53060 56028 54012 56084
rect 54068 56028 54078 56084
rect 12898 55916 12908 55972
rect 12964 55916 14140 55972
rect 14196 55916 17836 55972
rect 17892 55916 17902 55972
rect 18834 55916 18844 55972
rect 18900 55916 25228 55972
rect 25284 55916 25294 55972
rect 30930 55916 30940 55972
rect 30996 55916 32396 55972
rect 32452 55916 32462 55972
rect 34290 55916 34300 55972
rect 34356 55916 35308 55972
rect 35364 55916 36092 55972
rect 36148 55916 36158 55972
rect 19170 55804 19180 55860
rect 19236 55804 19246 55860
rect 21746 55804 21756 55860
rect 21812 55804 24556 55860
rect 24612 55804 24622 55860
rect 24770 55804 24780 55860
rect 24836 55804 28700 55860
rect 28756 55804 28766 55860
rect 19180 55748 19236 55804
rect 12786 55692 12796 55748
rect 12852 55692 18844 55748
rect 18900 55692 18910 55748
rect 19180 55692 29484 55748
rect 29540 55692 29550 55748
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 17826 55580 17836 55636
rect 17892 55580 19180 55636
rect 19236 55580 22540 55636
rect 22596 55580 22606 55636
rect 22754 55580 22764 55636
rect 22820 55580 27916 55636
rect 27972 55580 27982 55636
rect 18050 55468 18060 55524
rect 18116 55468 19068 55524
rect 19124 55468 19134 55524
rect 19730 55468 19740 55524
rect 19796 55468 23212 55524
rect 23268 55468 23278 55524
rect 28354 55468 28364 55524
rect 28420 55468 28430 55524
rect 31602 55468 31612 55524
rect 31668 55468 36540 55524
rect 36596 55468 36606 55524
rect 20748 55412 20804 55468
rect 28364 55412 28420 55468
rect 14130 55356 14140 55412
rect 14196 55356 15260 55412
rect 15316 55356 15326 55412
rect 20738 55356 20748 55412
rect 20804 55356 20814 55412
rect 22418 55356 22428 55412
rect 22484 55356 24332 55412
rect 24388 55356 24398 55412
rect 26114 55356 26124 55412
rect 26180 55356 26684 55412
rect 26740 55356 31724 55412
rect 31780 55356 31790 55412
rect 35970 55356 35980 55412
rect 36036 55356 37884 55412
rect 37940 55356 37950 55412
rect 14578 55244 14588 55300
rect 14644 55244 14654 55300
rect 14914 55244 14924 55300
rect 14980 55244 15036 55300
rect 15092 55244 15102 55300
rect 15362 55244 15372 55300
rect 15428 55244 15932 55300
rect 15988 55244 16604 55300
rect 16660 55244 18732 55300
rect 18788 55244 18798 55300
rect 20178 55244 20188 55300
rect 20244 55244 25340 55300
rect 25396 55244 25406 55300
rect 27570 55244 27580 55300
rect 27636 55244 28252 55300
rect 28308 55244 28318 55300
rect 38210 55244 38220 55300
rect 38276 55244 40348 55300
rect 40404 55244 41804 55300
rect 41860 55244 41870 55300
rect 42476 55244 43372 55300
rect 43428 55244 43438 55300
rect 14588 55188 14644 55244
rect 42476 55188 42532 55244
rect 14588 55132 15316 55188
rect 15586 55132 15596 55188
rect 15652 55132 17388 55188
rect 17444 55132 17454 55188
rect 22194 55132 22204 55188
rect 22260 55132 23548 55188
rect 23604 55132 23614 55188
rect 31042 55132 31052 55188
rect 31108 55132 32732 55188
rect 32788 55132 33180 55188
rect 33236 55132 34860 55188
rect 34916 55132 34926 55188
rect 36418 55132 36428 55188
rect 36484 55132 42476 55188
rect 42532 55132 42542 55188
rect 42690 55132 42700 55188
rect 42756 55132 43820 55188
rect 43876 55132 43886 55188
rect 4162 55020 4172 55076
rect 4228 55020 4732 55076
rect 4788 55020 12460 55076
rect 12516 55020 12526 55076
rect 15260 54964 15316 55132
rect 16482 55020 16492 55076
rect 16548 55020 16558 55076
rect 27570 55020 27580 55076
rect 27636 55020 29260 55076
rect 29316 55020 29820 55076
rect 29876 55020 29886 55076
rect 31686 55020 31724 55076
rect 31780 55020 34300 55076
rect 34356 55020 34366 55076
rect 36642 55020 36652 55076
rect 36708 55020 37324 55076
rect 37380 55020 37390 55076
rect 37986 55020 37996 55076
rect 38052 55020 38780 55076
rect 38836 55020 38846 55076
rect 42578 55020 42588 55076
rect 42644 55020 48188 55076
rect 48244 55020 48748 55076
rect 48804 55020 48814 55076
rect 16492 54964 16548 55020
rect 15260 54908 16548 54964
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 23762 54796 23772 54852
rect 23828 54796 24892 54852
rect 24948 54796 24958 54852
rect 26786 54796 26796 54852
rect 26852 54796 36988 54852
rect 37044 54796 37054 54852
rect 12002 54684 12012 54740
rect 12068 54684 12908 54740
rect 12964 54684 12974 54740
rect 22642 54684 22652 54740
rect 22708 54684 22718 54740
rect 26226 54684 26236 54740
rect 26292 54684 33628 54740
rect 33684 54684 33694 54740
rect 34738 54684 34748 54740
rect 34804 54684 38220 54740
rect 38276 54684 38286 54740
rect 45490 54684 45500 54740
rect 45556 54684 50764 54740
rect 50820 54684 51436 54740
rect 51492 54684 51884 54740
rect 51940 54684 51950 54740
rect 22652 54628 22708 54684
rect 12450 54572 12460 54628
rect 12516 54572 12526 54628
rect 14466 54572 14476 54628
rect 14532 54572 15372 54628
rect 15428 54572 15438 54628
rect 16706 54572 16716 54628
rect 16772 54572 21756 54628
rect 21812 54572 21822 54628
rect 22652 54572 30380 54628
rect 30436 54572 30446 54628
rect 37650 54572 37660 54628
rect 37716 54572 46396 54628
rect 46452 54572 46462 54628
rect 46946 54572 46956 54628
rect 47012 54572 49084 54628
rect 49140 54572 49150 54628
rect 0 54516 800 54544
rect 0 54460 1932 54516
rect 1988 54460 1998 54516
rect 0 54432 800 54460
rect 12460 54404 12516 54572
rect 46396 54516 46452 54572
rect 14242 54460 14252 54516
rect 14308 54460 14700 54516
rect 14756 54460 14766 54516
rect 17798 54460 17836 54516
rect 17892 54460 17902 54516
rect 18386 54460 18396 54516
rect 18452 54460 19740 54516
rect 19796 54460 19806 54516
rect 24546 54460 24556 54516
rect 24612 54460 26908 54516
rect 26964 54460 26974 54516
rect 28354 54460 28364 54516
rect 28420 54460 38220 54516
rect 38276 54460 38286 54516
rect 38612 54460 39788 54516
rect 39844 54460 42140 54516
rect 42196 54460 42206 54516
rect 42802 54460 42812 54516
rect 42868 54460 43708 54516
rect 43764 54460 43774 54516
rect 46396 54460 47628 54516
rect 47684 54460 47694 54516
rect 48290 54460 48300 54516
rect 48356 54460 48972 54516
rect 49028 54460 49038 54516
rect 49522 54460 49532 54516
rect 49588 54460 50652 54516
rect 50708 54460 54572 54516
rect 54628 54460 54638 54516
rect 11890 54348 11900 54404
rect 11956 54348 13580 54404
rect 13636 54348 15036 54404
rect 15092 54348 15102 54404
rect 16230 54348 16268 54404
rect 16324 54348 16334 54404
rect 23538 54348 23548 54404
rect 23604 54348 23884 54404
rect 23940 54348 23950 54404
rect 24658 54348 24668 54404
rect 24724 54348 26124 54404
rect 26180 54348 26190 54404
rect 30146 54348 30156 54404
rect 30212 54348 30604 54404
rect 30660 54348 31500 54404
rect 31556 54348 33964 54404
rect 34020 54348 34030 54404
rect 38612 54292 38668 54460
rect 38882 54348 38892 54404
rect 38948 54348 39564 54404
rect 39620 54348 39630 54404
rect 42690 54348 42700 54404
rect 42756 54348 44492 54404
rect 44548 54348 49196 54404
rect 49252 54348 49262 54404
rect 50866 54348 50876 54404
rect 50932 54348 53228 54404
rect 53284 54348 53294 54404
rect 17042 54236 17052 54292
rect 17108 54236 18172 54292
rect 18228 54236 18238 54292
rect 22082 54236 22092 54292
rect 22148 54236 24220 54292
rect 24276 54236 24286 54292
rect 28354 54236 28364 54292
rect 28420 54236 30268 54292
rect 30324 54236 30334 54292
rect 30594 54236 30604 54292
rect 30660 54236 30670 54292
rect 31826 54236 31836 54292
rect 31892 54236 38668 54292
rect 41906 54236 41916 54292
rect 41972 54236 44940 54292
rect 44996 54236 45006 54292
rect 47842 54236 47852 54292
rect 47908 54236 49868 54292
rect 49924 54236 49934 54292
rect 30604 54180 30660 54236
rect 6514 54124 6524 54180
rect 6580 54124 27580 54180
rect 27636 54124 27646 54180
rect 30370 54124 30380 54180
rect 30436 54124 30660 54180
rect 33618 54124 33628 54180
rect 33684 54124 34300 54180
rect 34356 54124 34366 54180
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 12898 54012 12908 54068
rect 12964 54012 15932 54068
rect 15988 54012 17052 54068
rect 17108 54012 17118 54068
rect 17378 54012 17388 54068
rect 17444 54012 19628 54068
rect 19684 54012 28140 54068
rect 28196 54012 28206 54068
rect 13122 53900 13132 53956
rect 13188 53900 15148 53956
rect 16482 53900 16492 53956
rect 16548 53900 18340 53956
rect 19394 53900 19404 53956
rect 19460 53900 21196 53956
rect 21252 53900 21262 53956
rect 21420 53900 29596 53956
rect 29652 53900 29820 53956
rect 29876 53900 29932 53956
rect 29988 53900 29998 53956
rect 33170 53900 33180 53956
rect 33236 53900 34076 53956
rect 34132 53900 34142 53956
rect 35410 53900 35420 53956
rect 35476 53900 37212 53956
rect 37268 53900 37278 53956
rect 39778 53900 39788 53956
rect 39844 53900 40684 53956
rect 40740 53900 42028 53956
rect 42084 53900 42094 53956
rect 46834 53900 46844 53956
rect 46900 53900 47516 53956
rect 47572 53900 48076 53956
rect 48132 53900 48142 53956
rect 15092 53844 15148 53900
rect 18284 53844 18340 53900
rect 21420 53844 21476 53900
rect 15092 53788 18060 53844
rect 18116 53788 18126 53844
rect 18284 53788 20412 53844
rect 20468 53788 21476 53844
rect 23090 53788 23100 53844
rect 23156 53788 23436 53844
rect 23492 53788 23502 53844
rect 28130 53788 28140 53844
rect 28196 53788 31164 53844
rect 31220 53788 31230 53844
rect 35186 53788 35196 53844
rect 35252 53788 36204 53844
rect 36260 53788 36764 53844
rect 36820 53788 36830 53844
rect 40002 53788 40012 53844
rect 40068 53788 40796 53844
rect 40852 53788 40862 53844
rect 46498 53788 46508 53844
rect 46564 53788 47068 53844
rect 47124 53788 47740 53844
rect 47796 53788 47806 53844
rect 15092 53676 15708 53732
rect 15764 53676 15774 53732
rect 23650 53676 23660 53732
rect 23716 53676 24108 53732
rect 24164 53676 24174 53732
rect 26002 53676 26012 53732
rect 26068 53676 26684 53732
rect 26740 53676 26750 53732
rect 30146 53676 30156 53732
rect 30212 53676 32956 53732
rect 33012 53676 33022 53732
rect 38994 53676 39004 53732
rect 39060 53676 42252 53732
rect 42308 53676 43260 53732
rect 43316 53676 43326 53732
rect 45826 53676 45836 53732
rect 45892 53676 47180 53732
rect 47236 53676 47246 53732
rect 51090 53676 51100 53732
rect 51156 53676 52780 53732
rect 52836 53676 52846 53732
rect 53890 53676 53900 53732
rect 53956 53676 55580 53732
rect 55636 53676 55646 53732
rect 13318 53564 13356 53620
rect 13412 53564 13422 53620
rect 15092 53508 15148 53676
rect 22418 53564 22428 53620
rect 22484 53564 22988 53620
rect 23044 53564 23054 53620
rect 26450 53564 26460 53620
rect 26516 53564 29148 53620
rect 29204 53564 29214 53620
rect 29586 53564 29596 53620
rect 29652 53564 32172 53620
rect 32228 53564 32238 53620
rect 33282 53564 33292 53620
rect 33348 53564 34524 53620
rect 34580 53564 34590 53620
rect 36082 53564 36092 53620
rect 36148 53564 36876 53620
rect 36932 53564 36942 53620
rect 40338 53564 40348 53620
rect 40404 53564 41356 53620
rect 41412 53564 41422 53620
rect 42466 53564 42476 53620
rect 42532 53564 43148 53620
rect 43204 53564 43214 53620
rect 47618 53564 47628 53620
rect 47684 53564 50092 53620
rect 50148 53564 50158 53620
rect 8306 53452 8316 53508
rect 8372 53396 8428 53508
rect 10658 53452 10668 53508
rect 10724 53452 14476 53508
rect 14532 53452 14812 53508
rect 14868 53452 15148 53508
rect 17154 53452 17164 53508
rect 17220 53452 18844 53508
rect 18900 53452 24668 53508
rect 24724 53452 24734 53508
rect 26562 53452 26572 53508
rect 26628 53452 26908 53508
rect 26964 53452 27860 53508
rect 28018 53452 28028 53508
rect 28084 53452 30940 53508
rect 30996 53452 31006 53508
rect 31154 53452 31164 53508
rect 31220 53452 31724 53508
rect 31780 53452 31790 53508
rect 33842 53452 33852 53508
rect 33908 53452 35980 53508
rect 36036 53452 36046 53508
rect 38994 53452 39004 53508
rect 39060 53452 39676 53508
rect 39732 53452 39742 53508
rect 27804 53396 27860 53452
rect 8372 53340 10892 53396
rect 10948 53340 10958 53396
rect 11890 53340 11900 53396
rect 11956 53340 17500 53396
rect 17556 53340 17566 53396
rect 23538 53340 23548 53396
rect 23604 53340 26908 53396
rect 27804 53340 28364 53396
rect 28420 53340 28430 53396
rect 29810 53340 29820 53396
rect 29876 53340 31612 53396
rect 31668 53340 31678 53396
rect 11900 53284 11956 53340
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 26852 53284 26908 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 9762 53228 9772 53284
rect 9828 53228 11956 53284
rect 13682 53228 13692 53284
rect 13748 53228 17836 53284
rect 17892 53228 17902 53284
rect 26852 53228 30604 53284
rect 30660 53228 30670 53284
rect 59200 53172 60000 53200
rect 13346 53116 13356 53172
rect 13412 53116 15484 53172
rect 15540 53116 15550 53172
rect 17490 53116 17500 53172
rect 17556 53116 17612 53172
rect 17668 53116 24332 53172
rect 24388 53116 24398 53172
rect 28018 53116 28028 53172
rect 28084 53116 29484 53172
rect 29540 53116 29550 53172
rect 31154 53116 31164 53172
rect 31220 53116 31948 53172
rect 32004 53116 32014 53172
rect 33590 53116 33628 53172
rect 33684 53116 34860 53172
rect 34916 53116 35420 53172
rect 35476 53116 35486 53172
rect 36978 53116 36988 53172
rect 37044 53116 37996 53172
rect 38052 53116 38444 53172
rect 38500 53116 39564 53172
rect 39620 53116 40124 53172
rect 40180 53116 40190 53172
rect 57250 53116 57260 53172
rect 57316 53116 60000 53172
rect 59200 53088 60000 53116
rect 13346 53004 13356 53060
rect 13412 53004 15148 53060
rect 19394 53004 19404 53060
rect 19460 53004 22540 53060
rect 22596 53004 24444 53060
rect 24500 53004 24510 53060
rect 24658 53004 24668 53060
rect 24724 53004 25116 53060
rect 25172 53004 29036 53060
rect 29092 53004 29102 53060
rect 30706 53004 30716 53060
rect 30772 53004 34972 53060
rect 35028 53004 38668 53060
rect 38882 53004 38892 53060
rect 38948 53004 39228 53060
rect 39284 53004 39452 53060
rect 39508 53004 40012 53060
rect 40068 53004 40078 53060
rect 50082 53004 50092 53060
rect 50148 53004 51548 53060
rect 51604 53004 51614 53060
rect 15092 52948 15148 53004
rect 38612 52948 38668 53004
rect 11330 52892 11340 52948
rect 11396 52892 12124 52948
rect 12180 52892 12190 52948
rect 12562 52892 12572 52948
rect 12628 52892 13916 52948
rect 13972 52892 14252 52948
rect 14308 52892 14318 52948
rect 15092 52892 21308 52948
rect 21364 52892 21374 52948
rect 27346 52892 27356 52948
rect 27412 52892 36428 52948
rect 36484 52892 36494 52948
rect 38612 52892 39004 52948
rect 39060 52892 39070 52948
rect 13766 52780 13804 52836
rect 13860 52780 13870 52836
rect 16370 52780 16380 52836
rect 16436 52780 17276 52836
rect 17332 52780 19572 52836
rect 19730 52780 19740 52836
rect 19796 52780 20188 52836
rect 20244 52780 21644 52836
rect 21700 52780 21710 52836
rect 23314 52780 23324 52836
rect 23380 52780 25564 52836
rect 25620 52780 25630 52836
rect 26562 52780 26572 52836
rect 26628 52780 28308 52836
rect 28914 52780 28924 52836
rect 28980 52780 36988 52836
rect 37044 52780 37054 52836
rect 19516 52724 19572 52780
rect 11778 52668 11788 52724
rect 11844 52668 12348 52724
rect 12404 52668 15148 52724
rect 16034 52668 16044 52724
rect 16100 52668 18620 52724
rect 18676 52668 18686 52724
rect 19516 52668 23660 52724
rect 23716 52668 23726 52724
rect 15092 52612 15148 52668
rect 28252 52612 28308 52780
rect 31826 52668 31836 52724
rect 31892 52668 33068 52724
rect 33124 52668 33134 52724
rect 34486 52668 34524 52724
rect 34580 52668 34590 52724
rect 15092 52556 17164 52612
rect 17220 52556 18284 52612
rect 18340 52556 18350 52612
rect 23650 52556 23660 52612
rect 23716 52556 24780 52612
rect 24836 52556 27580 52612
rect 27636 52556 27646 52612
rect 28242 52556 28252 52612
rect 28308 52556 28318 52612
rect 28578 52556 28588 52612
rect 28644 52556 32060 52612
rect 32116 52556 32126 52612
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 12338 52444 12348 52500
rect 12404 52444 17052 52500
rect 17108 52444 17118 52500
rect 20710 52444 20748 52500
rect 20804 52444 20814 52500
rect 21410 52444 21420 52500
rect 21476 52444 26460 52500
rect 26516 52444 26526 52500
rect 28018 52444 28028 52500
rect 28084 52444 28476 52500
rect 28532 52444 28542 52500
rect 32060 52388 32116 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 43260 52444 45612 52500
rect 45668 52444 45678 52500
rect 11106 52332 11116 52388
rect 11172 52332 12460 52388
rect 12516 52332 12526 52388
rect 18050 52332 18060 52388
rect 18116 52332 19068 52388
rect 19124 52332 26012 52388
rect 26068 52332 26078 52388
rect 26674 52332 26684 52388
rect 26740 52332 28644 52388
rect 32060 52332 35644 52388
rect 35700 52332 35710 52388
rect 37986 52332 37996 52388
rect 38052 52332 41244 52388
rect 41300 52332 41310 52388
rect 41682 52332 41692 52388
rect 41748 52332 42476 52388
rect 42532 52332 42542 52388
rect 8754 52220 8764 52276
rect 8820 52220 10780 52276
rect 10836 52220 10846 52276
rect 14326 52220 14364 52276
rect 14420 52220 14430 52276
rect 17602 52220 17612 52276
rect 17668 52220 19180 52276
rect 19236 52220 19246 52276
rect 19590 52220 19628 52276
rect 19684 52220 19694 52276
rect 20178 52220 20188 52276
rect 20244 52220 21420 52276
rect 21476 52220 21486 52276
rect 22978 52220 22988 52276
rect 23044 52220 26796 52276
rect 26852 52220 27916 52276
rect 27972 52220 27982 52276
rect 8530 52108 8540 52164
rect 8596 52108 9324 52164
rect 9380 52108 10332 52164
rect 10388 52108 10398 52164
rect 14018 52108 14028 52164
rect 14084 52108 16156 52164
rect 16212 52108 16222 52164
rect 20290 52108 20300 52164
rect 20356 52108 21084 52164
rect 21140 52108 21150 52164
rect 21634 52108 21644 52164
rect 21700 52108 22540 52164
rect 22596 52108 23660 52164
rect 23716 52108 23726 52164
rect 23986 52108 23996 52164
rect 24052 52108 25676 52164
rect 25732 52108 27132 52164
rect 27188 52108 27198 52164
rect 15446 51996 15484 52052
rect 15540 51996 15550 52052
rect 18274 51996 18284 52052
rect 18340 51996 26124 52052
rect 26180 51996 26190 52052
rect 28588 51940 28644 52332
rect 43260 52276 43316 52444
rect 43922 52332 43932 52388
rect 43988 52332 46172 52388
rect 46228 52332 46238 52388
rect 31826 52220 31836 52276
rect 31892 52220 39452 52276
rect 39508 52220 39518 52276
rect 41010 52220 41020 52276
rect 41076 52220 43260 52276
rect 43316 52220 43326 52276
rect 43474 52220 43484 52276
rect 43540 52220 44044 52276
rect 44100 52220 45164 52276
rect 45220 52220 45230 52276
rect 47394 52220 47404 52276
rect 47460 52220 48188 52276
rect 48244 52220 49084 52276
rect 49140 52220 50204 52276
rect 50260 52220 50270 52276
rect 30790 52108 30828 52164
rect 30884 52108 30894 52164
rect 34850 52108 34860 52164
rect 34916 52108 35420 52164
rect 35476 52108 35486 52164
rect 40226 52108 40236 52164
rect 40292 52108 41132 52164
rect 41188 52108 41198 52164
rect 43586 52108 43596 52164
rect 43652 52108 44828 52164
rect 44884 52108 44894 52164
rect 48850 52108 48860 52164
rect 48916 52108 50428 52164
rect 50484 52108 50988 52164
rect 51044 52108 51054 52164
rect 43250 51996 43260 52052
rect 43316 51996 43484 52052
rect 43540 51996 43550 52052
rect 50306 51996 50316 52052
rect 50372 51996 51212 52052
rect 51268 51996 51278 52052
rect 15092 51884 18060 51940
rect 18116 51884 20468 51940
rect 20598 51884 20636 51940
rect 20692 51884 20702 51940
rect 20850 51884 20860 51940
rect 20916 51884 20954 51940
rect 28588 51884 29260 51940
rect 29316 51884 29708 51940
rect 29764 51884 29774 51940
rect 30370 51884 30380 51940
rect 30436 51884 31388 51940
rect 31444 51884 31454 51940
rect 37538 51884 37548 51940
rect 37604 51884 38444 51940
rect 38500 51884 38510 51940
rect 39666 51884 39676 51940
rect 39732 51884 42700 51940
rect 42756 51884 42766 51940
rect 15092 51716 15148 51884
rect 20412 51828 20468 51884
rect 20412 51772 21196 51828
rect 21252 51772 21262 51828
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 11442 51660 11452 51716
rect 11508 51660 12348 51716
rect 12404 51660 15148 51716
rect 24098 51660 24108 51716
rect 24164 51660 29036 51716
rect 29092 51660 29102 51716
rect 29932 51660 42476 51716
rect 42532 51660 42542 51716
rect 29932 51604 29988 51660
rect 18722 51548 18732 51604
rect 18788 51548 21868 51604
rect 21924 51548 25228 51604
rect 25284 51548 25294 51604
rect 29922 51548 29932 51604
rect 29988 51548 29998 51604
rect 30146 51548 30156 51604
rect 30212 51548 30604 51604
rect 30660 51548 30670 51604
rect 32946 51548 32956 51604
rect 33012 51548 33740 51604
rect 33796 51548 35196 51604
rect 35252 51548 35262 51604
rect 40898 51548 40908 51604
rect 40964 51548 47068 51604
rect 47124 51548 47134 51604
rect 9986 51436 9996 51492
rect 10052 51436 15260 51492
rect 15316 51436 15484 51492
rect 15540 51436 16156 51492
rect 16212 51436 16222 51492
rect 18050 51436 18060 51492
rect 18116 51436 20636 51492
rect 20692 51436 20702 51492
rect 21746 51436 21756 51492
rect 21812 51436 22316 51492
rect 22372 51436 31332 51492
rect 34850 51436 34860 51492
rect 34916 51436 37324 51492
rect 37380 51436 37390 51492
rect 38098 51436 38108 51492
rect 38164 51436 48636 51492
rect 48692 51436 48702 51492
rect 31276 51380 31332 51436
rect 8194 51324 8204 51380
rect 8260 51324 9548 51380
rect 9604 51324 11116 51380
rect 11172 51324 12684 51380
rect 12740 51324 12750 51380
rect 13234 51324 13244 51380
rect 13300 51324 14140 51380
rect 14196 51324 17724 51380
rect 17780 51324 17790 51380
rect 17938 51324 17948 51380
rect 18004 51324 18732 51380
rect 18788 51324 19180 51380
rect 19236 51324 19246 51380
rect 20178 51324 20188 51380
rect 20244 51324 20300 51380
rect 20356 51324 20366 51380
rect 20710 51324 20748 51380
rect 20804 51324 20814 51380
rect 21186 51324 21196 51380
rect 21252 51324 22708 51380
rect 22838 51324 22876 51380
rect 22932 51324 22942 51380
rect 23538 51324 23548 51380
rect 23604 51324 23614 51380
rect 24210 51324 24220 51380
rect 24276 51324 24668 51380
rect 24724 51324 24734 51380
rect 25218 51324 25228 51380
rect 25284 51324 26124 51380
rect 26180 51324 26190 51380
rect 27094 51324 27132 51380
rect 27188 51324 27198 51380
rect 31266 51324 31276 51380
rect 31332 51324 31342 51380
rect 22652 51268 22708 51324
rect 23548 51268 23604 51324
rect 16370 51212 16380 51268
rect 16436 51212 18844 51268
rect 18900 51212 18910 51268
rect 20402 51212 20412 51268
rect 20468 51212 21644 51268
rect 21700 51212 21710 51268
rect 22652 51212 24108 51268
rect 24164 51212 24174 51268
rect 26562 51212 26572 51268
rect 26628 51212 27804 51268
rect 27860 51212 27870 51268
rect 41682 51212 41692 51268
rect 41748 51212 45836 51268
rect 45892 51212 45902 51268
rect 46498 51212 46508 51268
rect 46564 51212 46956 51268
rect 47012 51212 47516 51268
rect 47572 51212 47582 51268
rect 0 51156 800 51184
rect 0 51100 1708 51156
rect 1764 51100 1774 51156
rect 16818 51100 16828 51156
rect 16884 51100 18732 51156
rect 18788 51100 18798 51156
rect 20066 51100 20076 51156
rect 20132 51100 20142 51156
rect 22530 51100 22540 51156
rect 22596 51100 23548 51156
rect 23604 51100 23614 51156
rect 26852 51100 29820 51156
rect 29876 51100 29886 51156
rect 31378 51100 31388 51156
rect 31444 51100 32060 51156
rect 32116 51100 33292 51156
rect 33348 51100 33358 51156
rect 43026 51100 43036 51156
rect 43092 51100 43708 51156
rect 43764 51100 43774 51156
rect 0 51072 800 51100
rect 20076 51044 20132 51100
rect 26852 51044 26908 51100
rect 20076 50988 26908 51044
rect 27244 50988 29372 51044
rect 29428 50988 31612 51044
rect 31668 50988 32284 51044
rect 32340 50988 33180 51044
rect 33236 50988 33246 51044
rect 37090 50988 37100 51044
rect 37156 50988 37772 51044
rect 37828 50988 37838 51044
rect 42690 50988 42700 51044
rect 42756 50988 43484 51044
rect 43540 50988 43550 51044
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 27244 50932 27300 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 16706 50876 16716 50932
rect 16772 50876 20188 50932
rect 20244 50876 20254 50932
rect 20626 50876 20636 50932
rect 20692 50876 24892 50932
rect 24948 50876 26404 50932
rect 26674 50876 26684 50932
rect 26740 50876 27300 50932
rect 30034 50876 30044 50932
rect 30100 50876 34188 50932
rect 34244 50876 34254 50932
rect 36978 50876 36988 50932
rect 37044 50876 38668 50932
rect 26348 50820 26404 50876
rect 13570 50764 13580 50820
rect 13636 50764 16940 50820
rect 16996 50764 17006 50820
rect 18508 50764 23884 50820
rect 23940 50764 26124 50820
rect 26180 50764 26190 50820
rect 26348 50764 27916 50820
rect 27972 50764 27982 50820
rect 30146 50764 30156 50820
rect 30212 50764 30716 50820
rect 30772 50764 30782 50820
rect 31154 50764 31164 50820
rect 31220 50764 38108 50820
rect 38164 50764 38174 50820
rect 18508 50708 18564 50764
rect 38612 50708 38668 50876
rect 9538 50652 9548 50708
rect 9604 50652 14252 50708
rect 14308 50652 14318 50708
rect 15026 50652 15036 50708
rect 15092 50652 18564 50708
rect 18722 50652 18732 50708
rect 18788 50652 21196 50708
rect 21252 50652 21262 50708
rect 23762 50652 23772 50708
rect 23828 50652 24892 50708
rect 24948 50652 25788 50708
rect 25844 50652 25854 50708
rect 26852 50652 32284 50708
rect 32340 50652 32350 50708
rect 35186 50652 35196 50708
rect 35252 50652 37436 50708
rect 37492 50652 38332 50708
rect 38388 50652 38398 50708
rect 38612 50652 39564 50708
rect 39620 50652 39630 50708
rect 47506 50652 47516 50708
rect 47572 50652 48076 50708
rect 48132 50652 48142 50708
rect 49634 50652 49644 50708
rect 49700 50652 50652 50708
rect 50708 50652 51212 50708
rect 51268 50652 51278 50708
rect 51986 50652 51996 50708
rect 52052 50652 52332 50708
rect 52388 50652 52668 50708
rect 52724 50652 52734 50708
rect 14252 50596 14308 50652
rect 26852 50596 26908 50652
rect 12226 50540 12236 50596
rect 12292 50540 13692 50596
rect 13748 50540 13758 50596
rect 14252 50540 15596 50596
rect 15652 50540 15662 50596
rect 17490 50540 17500 50596
rect 17556 50540 18060 50596
rect 18116 50540 18126 50596
rect 18610 50540 18620 50596
rect 18676 50540 19628 50596
rect 19684 50540 22204 50596
rect 22260 50540 22270 50596
rect 23986 50540 23996 50596
rect 24052 50540 24062 50596
rect 24294 50540 24332 50596
rect 24388 50540 24398 50596
rect 25554 50540 25564 50596
rect 25620 50540 26908 50596
rect 27346 50540 27356 50596
rect 27412 50540 27422 50596
rect 30006 50540 30044 50596
rect 30100 50540 30110 50596
rect 30258 50540 30268 50596
rect 30324 50540 31052 50596
rect 31108 50540 33740 50596
rect 33796 50540 33806 50596
rect 34178 50540 34188 50596
rect 34244 50540 36372 50596
rect 37986 50540 37996 50596
rect 38052 50540 43260 50596
rect 43316 50540 43326 50596
rect 45602 50540 45612 50596
rect 45668 50540 46060 50596
rect 46116 50540 46284 50596
rect 46340 50540 46350 50596
rect 47282 50540 47292 50596
rect 47348 50540 49084 50596
rect 49140 50540 50092 50596
rect 50148 50540 50158 50596
rect 23996 50484 24052 50540
rect 27356 50484 27412 50540
rect 36316 50484 36372 50540
rect 59200 50484 60000 50512
rect 10098 50428 10108 50484
rect 10164 50428 10444 50484
rect 10500 50428 16380 50484
rect 16436 50428 16446 50484
rect 20738 50428 20748 50484
rect 20804 50428 21084 50484
rect 21140 50428 24052 50484
rect 24434 50428 24444 50484
rect 24500 50428 27412 50484
rect 29148 50428 30604 50484
rect 30660 50428 30670 50484
rect 31350 50428 31388 50484
rect 31444 50428 31454 50484
rect 32162 50428 32172 50484
rect 32228 50428 32732 50484
rect 32788 50428 32798 50484
rect 36306 50428 36316 50484
rect 36372 50428 38780 50484
rect 38836 50428 38846 50484
rect 44258 50428 44268 50484
rect 44324 50428 45948 50484
rect 46004 50428 46732 50484
rect 46788 50428 46798 50484
rect 46946 50428 46956 50484
rect 47012 50428 48860 50484
rect 48916 50428 49420 50484
rect 49476 50428 49486 50484
rect 50194 50428 50204 50484
rect 50260 50428 50764 50484
rect 50820 50428 50830 50484
rect 57820 50428 60000 50484
rect 21868 50372 21924 50428
rect 29148 50372 29204 50428
rect 57820 50372 57876 50428
rect 59200 50400 60000 50428
rect 18722 50316 18732 50372
rect 18788 50316 19628 50372
rect 19684 50316 19694 50372
rect 19954 50316 19964 50372
rect 20020 50316 21420 50372
rect 21476 50316 21486 50372
rect 21634 50316 21644 50372
rect 21700 50316 21924 50372
rect 22978 50316 22988 50372
rect 23044 50316 26236 50372
rect 26292 50316 26302 50372
rect 26786 50316 26796 50372
rect 26852 50316 27132 50372
rect 27188 50316 27198 50372
rect 27346 50316 27356 50372
rect 27412 50316 29204 50372
rect 29362 50316 29372 50372
rect 29428 50316 32620 50372
rect 32676 50316 32686 50372
rect 32834 50316 32844 50372
rect 32900 50316 33516 50372
rect 33572 50316 33582 50372
rect 42802 50316 42812 50372
rect 42868 50316 43596 50372
rect 43652 50316 43662 50372
rect 52882 50316 52892 50372
rect 52948 50316 54348 50372
rect 54404 50316 54414 50372
rect 57810 50316 57820 50372
rect 57876 50316 57886 50372
rect 13010 50204 13020 50260
rect 13076 50204 16828 50260
rect 16884 50204 16894 50260
rect 20514 50204 20524 50260
rect 20580 50204 20860 50260
rect 20916 50204 20926 50260
rect 25890 50204 25900 50260
rect 25956 50204 30716 50260
rect 30772 50204 30782 50260
rect 40450 50204 40460 50260
rect 40516 50204 41020 50260
rect 41076 50204 42140 50260
rect 42196 50204 43372 50260
rect 43428 50204 43438 50260
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 11666 50092 11676 50148
rect 11732 50092 16604 50148
rect 16660 50092 16670 50148
rect 18806 50092 18844 50148
rect 18900 50092 18910 50148
rect 20188 50092 25676 50148
rect 25732 50092 25742 50148
rect 26002 50092 26012 50148
rect 26068 50092 26460 50148
rect 26516 50092 26526 50148
rect 26898 50092 26908 50148
rect 26964 50092 27244 50148
rect 27300 50092 27310 50148
rect 27458 50092 27468 50148
rect 27524 50092 29596 50148
rect 29652 50092 29662 50148
rect 31714 50092 31724 50148
rect 31780 50092 32508 50148
rect 32564 50092 32574 50148
rect 20188 50036 20244 50092
rect 13794 49980 13804 50036
rect 13860 49980 15260 50036
rect 15316 49980 15326 50036
rect 17378 49980 17388 50036
rect 17444 49980 18732 50036
rect 18788 49980 20244 50036
rect 22978 49980 22988 50036
rect 23044 49980 38444 50036
rect 38500 49980 38510 50036
rect 40562 49980 40572 50036
rect 40628 49980 41468 50036
rect 41524 49980 44380 50036
rect 44436 49980 44446 50036
rect 16818 49868 16828 49924
rect 16884 49868 20188 49924
rect 20244 49868 21084 49924
rect 21140 49868 21150 49924
rect 23090 49868 23100 49924
rect 23156 49868 23660 49924
rect 23716 49868 23726 49924
rect 24658 49868 24668 49924
rect 24724 49868 25564 49924
rect 25620 49868 25630 49924
rect 26562 49868 26572 49924
rect 26628 49868 30380 49924
rect 30436 49868 30446 49924
rect 30604 49868 31276 49924
rect 31332 49868 32396 49924
rect 32452 49868 32462 49924
rect 43362 49868 43372 49924
rect 43428 49868 45276 49924
rect 45332 49868 45342 49924
rect 54226 49868 54236 49924
rect 54292 49868 54908 49924
rect 54964 49868 54974 49924
rect 30604 49812 30660 49868
rect 59200 49812 60000 49840
rect 8306 49756 8316 49812
rect 8372 49756 8876 49812
rect 8932 49756 9548 49812
rect 9604 49756 9614 49812
rect 17378 49756 17388 49812
rect 17444 49756 19292 49812
rect 19348 49756 19358 49812
rect 20402 49756 20412 49812
rect 20468 49756 22764 49812
rect 22820 49756 22830 49812
rect 26786 49756 26796 49812
rect 26852 49756 26862 49812
rect 27206 49756 27244 49812
rect 27300 49756 28028 49812
rect 28084 49756 28094 49812
rect 28242 49756 28252 49812
rect 28308 49756 29372 49812
rect 29428 49756 30660 49812
rect 30818 49756 30828 49812
rect 30884 49756 31388 49812
rect 31444 49756 31454 49812
rect 35410 49756 35420 49812
rect 35476 49756 36316 49812
rect 36372 49756 36652 49812
rect 36708 49756 36718 49812
rect 40226 49756 40236 49812
rect 40292 49756 46844 49812
rect 46900 49756 46910 49812
rect 51762 49756 51772 49812
rect 51828 49756 53004 49812
rect 53060 49756 53900 49812
rect 53956 49756 53966 49812
rect 57922 49756 57932 49812
rect 57988 49756 60000 49812
rect 26796 49700 26852 49756
rect 59200 49728 60000 49756
rect 16258 49644 16268 49700
rect 16324 49644 18284 49700
rect 18340 49644 18350 49700
rect 19954 49644 19964 49700
rect 20020 49644 22092 49700
rect 22148 49644 22158 49700
rect 22316 49644 26852 49700
rect 27766 49644 27804 49700
rect 27860 49644 27870 49700
rect 29474 49644 29484 49700
rect 29540 49644 34972 49700
rect 35028 49644 35038 49700
rect 22316 49588 22372 49644
rect 15250 49532 15260 49588
rect 15316 49532 21308 49588
rect 21364 49532 21374 49588
rect 21634 49532 21644 49588
rect 21700 49532 22372 49588
rect 26786 49532 26796 49588
rect 26852 49532 36876 49588
rect 36932 49532 36942 49588
rect 10434 49420 10444 49476
rect 10500 49420 12012 49476
rect 12068 49420 19852 49476
rect 19908 49420 23324 49476
rect 23380 49420 23390 49476
rect 26002 49420 26012 49476
rect 26068 49420 28364 49476
rect 28420 49420 28430 49476
rect 28914 49420 28924 49476
rect 28980 49420 30156 49476
rect 30212 49420 30222 49476
rect 30818 49420 30828 49476
rect 30884 49420 30940 49476
rect 30996 49420 31006 49476
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 11442 49308 11452 49364
rect 11508 49308 19180 49364
rect 19236 49308 19246 49364
rect 24098 49308 24108 49364
rect 24164 49308 24556 49364
rect 24612 49308 26908 49364
rect 26964 49308 31164 49364
rect 31220 49308 31230 49364
rect 10546 49196 10556 49252
rect 10612 49196 11116 49252
rect 11172 49196 12572 49252
rect 12628 49196 13580 49252
rect 13636 49196 13646 49252
rect 14690 49196 14700 49252
rect 14756 49196 21028 49252
rect 27570 49196 27580 49252
rect 27636 49196 28252 49252
rect 28308 49196 28318 49252
rect 40338 49196 40348 49252
rect 40404 49196 44268 49252
rect 44324 49196 44334 49252
rect 20178 49084 20188 49140
rect 20244 49084 20524 49140
rect 20580 49084 20590 49140
rect 20972 49028 21028 49196
rect 24220 49084 30828 49140
rect 30884 49084 30894 49140
rect 36418 49084 36428 49140
rect 36484 49084 37324 49140
rect 37380 49084 37390 49140
rect 37986 49084 37996 49140
rect 38052 49084 38444 49140
rect 38500 49084 38510 49140
rect 45378 49084 45388 49140
rect 45444 49084 46228 49140
rect 53106 49084 53116 49140
rect 53172 49084 53900 49140
rect 53956 49084 53966 49140
rect 24220 49028 24276 49084
rect 46172 49028 46228 49084
rect 11554 48972 11564 49028
rect 11620 48972 13580 49028
rect 13636 48972 13646 49028
rect 14578 48972 14588 49028
rect 14644 48972 15708 49028
rect 15764 48972 15774 49028
rect 16818 48972 16828 49028
rect 16884 48972 17500 49028
rect 17556 48972 17566 49028
rect 19954 48972 19964 49028
rect 20020 48972 20636 49028
rect 20692 48972 20702 49028
rect 20962 48972 20972 49028
rect 21028 48972 21308 49028
rect 21364 48972 21374 49028
rect 23314 48972 23324 49028
rect 23380 48972 24220 49028
rect 24276 48972 24286 49028
rect 25452 48972 26012 49028
rect 26068 48972 26078 49028
rect 26562 48972 26572 49028
rect 26628 48972 27804 49028
rect 27860 48972 27870 49028
rect 28326 48972 28364 49028
rect 28420 48972 28430 49028
rect 28578 48972 28588 49028
rect 28644 48972 29260 49028
rect 29316 48972 29326 49028
rect 30706 48972 30716 49028
rect 30772 48972 31948 49028
rect 32004 48972 33404 49028
rect 33460 48972 34412 49028
rect 34468 48972 34478 49028
rect 37884 48972 38668 49028
rect 39554 48972 39564 49028
rect 39620 48972 40908 49028
rect 40964 48972 40974 49028
rect 43810 48972 43820 49028
rect 43876 48972 45612 49028
rect 45668 48972 45678 49028
rect 46162 48972 46172 49028
rect 46228 48972 47180 49028
rect 47236 48972 47246 49028
rect 53666 48972 53676 49028
rect 53732 48972 54236 49028
rect 54292 48972 54302 49028
rect 25452 48916 25508 48972
rect 37884 48916 37940 48972
rect 38612 48916 38668 48972
rect 15810 48860 15820 48916
rect 15876 48860 16380 48916
rect 16436 48860 17724 48916
rect 17780 48860 18732 48916
rect 18788 48860 19628 48916
rect 19684 48860 19694 48916
rect 22540 48860 25508 48916
rect 25666 48860 25676 48916
rect 25732 48860 26908 48916
rect 27346 48860 27356 48916
rect 27412 48860 28868 48916
rect 37874 48860 37884 48916
rect 37940 48860 37950 48916
rect 38322 48860 38332 48916
rect 38388 48860 38398 48916
rect 38612 48860 39900 48916
rect 39956 48860 39966 48916
rect 43586 48860 43596 48916
rect 43652 48860 45836 48916
rect 45892 48860 45902 48916
rect 22540 48804 22596 48860
rect 26852 48804 26908 48860
rect 28812 48804 28868 48860
rect 38332 48804 38388 48860
rect 4274 48748 4284 48804
rect 4340 48748 4732 48804
rect 4788 48748 5628 48804
rect 5684 48748 5694 48804
rect 7858 48748 7868 48804
rect 7924 48748 8764 48804
rect 8820 48748 9548 48804
rect 9604 48748 9614 48804
rect 11106 48748 11116 48804
rect 11172 48748 12236 48804
rect 12292 48748 12302 48804
rect 16594 48748 16604 48804
rect 16660 48748 18508 48804
rect 18564 48748 22596 48804
rect 22754 48748 22764 48804
rect 22820 48748 24332 48804
rect 24388 48748 24398 48804
rect 25890 48748 25900 48804
rect 25956 48748 26684 48804
rect 26740 48748 26750 48804
rect 26852 48748 28028 48804
rect 28084 48748 28476 48804
rect 28532 48748 28542 48804
rect 28802 48748 28812 48804
rect 28868 48748 28878 48804
rect 29026 48748 29036 48804
rect 29092 48748 29820 48804
rect 29876 48748 30268 48804
rect 30324 48748 30334 48804
rect 31602 48748 31612 48804
rect 31668 48748 32396 48804
rect 32452 48748 32462 48804
rect 38332 48748 40460 48804
rect 40516 48748 40526 48804
rect 51986 48748 51996 48804
rect 52052 48748 52780 48804
rect 52836 48748 52846 48804
rect 16706 48636 16716 48692
rect 16772 48636 17724 48692
rect 17780 48636 17790 48692
rect 20262 48636 20300 48692
rect 20356 48636 20366 48692
rect 22866 48636 22876 48692
rect 22932 48636 29260 48692
rect 29316 48636 29326 48692
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 9874 48524 9884 48580
rect 9940 48524 12348 48580
rect 12404 48524 12414 48580
rect 27794 48524 27804 48580
rect 27860 48524 28252 48580
rect 28308 48524 28318 48580
rect 0 48468 800 48496
rect 0 48412 1932 48468
rect 1988 48412 1998 48468
rect 8082 48412 8092 48468
rect 8148 48412 10892 48468
rect 10948 48412 13468 48468
rect 13524 48412 13534 48468
rect 15362 48412 15372 48468
rect 15428 48412 24220 48468
rect 24276 48412 26572 48468
rect 26628 48412 26638 48468
rect 26786 48412 26796 48468
rect 26852 48412 27244 48468
rect 27300 48412 27310 48468
rect 28252 48412 29596 48468
rect 29652 48412 29662 48468
rect 29810 48412 29820 48468
rect 29876 48412 30268 48468
rect 30324 48412 30334 48468
rect 38210 48412 38220 48468
rect 38276 48412 38556 48468
rect 38612 48412 39004 48468
rect 39060 48412 39070 48468
rect 0 48384 800 48412
rect 28252 48356 28308 48412
rect 10658 48300 10668 48356
rect 10724 48300 12460 48356
rect 12516 48300 14476 48356
rect 14532 48300 14542 48356
rect 16818 48300 16828 48356
rect 16884 48300 17276 48356
rect 17332 48300 17342 48356
rect 24658 48300 24668 48356
rect 24724 48300 27468 48356
rect 27524 48300 27534 48356
rect 28018 48300 28028 48356
rect 28084 48300 28308 48356
rect 28364 48300 31052 48356
rect 31108 48300 31948 48356
rect 32004 48300 32014 48356
rect 48402 48300 48412 48356
rect 48468 48300 49420 48356
rect 49476 48300 49486 48356
rect 12338 48188 12348 48244
rect 12404 48188 15596 48244
rect 15652 48188 15662 48244
rect 18722 48188 18732 48244
rect 18788 48188 20076 48244
rect 20132 48188 21756 48244
rect 21812 48188 21822 48244
rect 25554 48188 25564 48244
rect 25620 48188 27244 48244
rect 27300 48188 27310 48244
rect 27654 48188 27692 48244
rect 27748 48188 27758 48244
rect 28364 48132 28420 48300
rect 29362 48188 29372 48244
rect 29428 48188 30268 48244
rect 30324 48188 30334 48244
rect 32946 48188 32956 48244
rect 33012 48188 34524 48244
rect 34580 48188 34590 48244
rect 44930 48188 44940 48244
rect 44996 48188 45612 48244
rect 45668 48188 46060 48244
rect 46116 48188 46126 48244
rect 47954 48188 47964 48244
rect 48020 48188 48972 48244
rect 49028 48188 50428 48244
rect 50484 48188 50494 48244
rect 52434 48188 52444 48244
rect 52500 48188 53228 48244
rect 53284 48188 53294 48244
rect 14802 48076 14812 48132
rect 14868 48076 20188 48132
rect 20244 48076 20254 48132
rect 21858 48076 21868 48132
rect 21924 48076 23100 48132
rect 23156 48076 23166 48132
rect 24098 48076 24108 48132
rect 24164 48076 28420 48132
rect 28578 48076 28588 48132
rect 28644 48076 31052 48132
rect 31108 48076 31118 48132
rect 32050 48076 32060 48132
rect 32116 48076 32844 48132
rect 32900 48076 32910 48132
rect 37090 48076 37100 48132
rect 37156 48076 37660 48132
rect 37716 48076 39452 48132
rect 39508 48076 39518 48132
rect 46274 48076 46284 48132
rect 46340 48076 46732 48132
rect 46788 48076 47740 48132
rect 47796 48076 47806 48132
rect 1922 47964 1932 48020
rect 1988 47964 1998 48020
rect 18694 47964 18732 48020
rect 18788 47964 18798 48020
rect 20626 47964 20636 48020
rect 20692 47964 21420 48020
rect 21476 47964 21486 48020
rect 25340 47964 25788 48020
rect 25844 47964 26572 48020
rect 26628 47964 26638 48020
rect 27542 47964 27580 48020
rect 27636 47964 27646 48020
rect 0 47796 800 47824
rect 1932 47796 1988 47964
rect 25340 47908 25396 47964
rect 28588 47908 28644 48076
rect 38108 48020 38164 48076
rect 38098 47964 38108 48020
rect 38164 47964 38174 48020
rect 38658 47964 38668 48020
rect 38724 47964 40348 48020
rect 40404 47964 40796 48020
rect 40852 47964 40862 48020
rect 46834 47964 46844 48020
rect 46900 47964 47404 48020
rect 47460 47964 47852 48020
rect 47908 47964 48860 48020
rect 48916 47964 48926 48020
rect 52658 47964 52668 48020
rect 52724 47964 53004 48020
rect 53060 47964 53070 48020
rect 16034 47852 16044 47908
rect 16100 47852 17948 47908
rect 18004 47852 25340 47908
rect 25396 47852 25406 47908
rect 25666 47852 25676 47908
rect 25732 47852 26796 47908
rect 26852 47852 28644 47908
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 0 47740 1988 47796
rect 11442 47740 11452 47796
rect 11508 47740 11518 47796
rect 18274 47740 18284 47796
rect 18340 47740 26684 47796
rect 26740 47740 26750 47796
rect 26852 47740 32844 47796
rect 32900 47740 33516 47796
rect 33572 47740 33582 47796
rect 0 47712 800 47740
rect 11452 47684 11508 47740
rect 11452 47628 11676 47684
rect 11732 47628 11742 47684
rect 16146 47628 16156 47684
rect 16212 47628 19012 47684
rect 19506 47628 19516 47684
rect 19572 47628 19852 47684
rect 19908 47628 20300 47684
rect 20356 47628 21644 47684
rect 21700 47628 21710 47684
rect 22306 47628 22316 47684
rect 22372 47628 25676 47684
rect 25732 47628 25742 47684
rect 18956 47572 19012 47628
rect 26852 47572 26908 47740
rect 27682 47628 27692 47684
rect 27748 47628 28364 47684
rect 28420 47628 29708 47684
rect 29764 47628 29774 47684
rect 30482 47628 30492 47684
rect 30548 47628 31164 47684
rect 31220 47628 31230 47684
rect 31714 47628 31724 47684
rect 31780 47628 35756 47684
rect 35812 47628 35980 47684
rect 36036 47628 36046 47684
rect 46162 47628 46172 47684
rect 46228 47628 47404 47684
rect 47460 47628 49532 47684
rect 49588 47628 50764 47684
rect 50820 47628 50830 47684
rect 11442 47516 11452 47572
rect 11508 47516 11788 47572
rect 11844 47516 11854 47572
rect 17042 47516 17052 47572
rect 17108 47516 18620 47572
rect 18676 47516 18686 47572
rect 18946 47516 18956 47572
rect 19012 47516 19022 47572
rect 20738 47516 20748 47572
rect 20804 47516 24108 47572
rect 24164 47516 24174 47572
rect 24658 47516 24668 47572
rect 24724 47516 26908 47572
rect 27234 47516 27244 47572
rect 27300 47516 29428 47572
rect 29586 47516 29596 47572
rect 29652 47516 31388 47572
rect 31444 47516 31454 47572
rect 33730 47516 33740 47572
rect 33796 47516 35308 47572
rect 35364 47516 35374 47572
rect 39330 47516 39340 47572
rect 39396 47516 40236 47572
rect 40292 47516 40302 47572
rect 29372 47460 29428 47516
rect 13122 47404 13132 47460
rect 13188 47404 15820 47460
rect 15876 47404 15886 47460
rect 16818 47404 16828 47460
rect 16884 47404 17388 47460
rect 17444 47404 17454 47460
rect 17714 47404 17724 47460
rect 17780 47404 22764 47460
rect 22820 47404 22830 47460
rect 22978 47404 22988 47460
rect 23044 47404 23772 47460
rect 23828 47404 23838 47460
rect 25218 47404 25228 47460
rect 25284 47404 26012 47460
rect 26068 47404 26078 47460
rect 26852 47404 28364 47460
rect 28420 47404 28430 47460
rect 29372 47404 33628 47460
rect 33684 47404 33694 47460
rect 37202 47404 37212 47460
rect 37268 47404 37436 47460
rect 37492 47404 38220 47460
rect 38276 47404 38286 47460
rect 45938 47404 45948 47460
rect 46004 47404 47180 47460
rect 47236 47404 48972 47460
rect 49028 47404 50204 47460
rect 50260 47404 50270 47460
rect 52098 47404 52108 47460
rect 52164 47404 52892 47460
rect 52948 47404 52958 47460
rect 26852 47348 26908 47404
rect 4274 47292 4284 47348
rect 4340 47292 7308 47348
rect 7364 47292 7374 47348
rect 14466 47292 14476 47348
rect 14532 47292 18284 47348
rect 18340 47292 19404 47348
rect 19460 47292 19470 47348
rect 23090 47292 23100 47348
rect 23156 47292 25452 47348
rect 25508 47292 26348 47348
rect 26404 47292 26908 47348
rect 28018 47292 28028 47348
rect 28084 47292 28094 47348
rect 29670 47292 29708 47348
rect 29764 47292 29774 47348
rect 30370 47292 30380 47348
rect 30436 47292 31724 47348
rect 31780 47292 32396 47348
rect 32452 47292 32462 47348
rect 34178 47292 34188 47348
rect 34244 47292 35868 47348
rect 35924 47292 35934 47348
rect 28028 47236 28084 47292
rect 8642 47180 8652 47236
rect 8708 47180 8876 47236
rect 8932 47180 9996 47236
rect 10052 47180 10062 47236
rect 16370 47180 16380 47236
rect 16436 47180 20412 47236
rect 20468 47180 20478 47236
rect 20738 47180 20748 47236
rect 20804 47180 28084 47236
rect 28466 47180 28476 47236
rect 28532 47180 32060 47236
rect 32116 47180 32126 47236
rect 51762 47180 51772 47236
rect 51828 47180 52220 47236
rect 52276 47180 52286 47236
rect 59200 47124 60000 47152
rect 11442 47068 11452 47124
rect 11508 47068 11732 47124
rect 11676 47012 11732 47068
rect 15092 47068 15484 47124
rect 15540 47068 18060 47124
rect 18116 47068 18126 47124
rect 18806 47068 18844 47124
rect 18900 47068 18910 47124
rect 20962 47068 20972 47124
rect 21028 47068 22540 47124
rect 22596 47068 23212 47124
rect 23268 47068 23278 47124
rect 27906 47068 27916 47124
rect 27972 47068 28252 47124
rect 28308 47068 29148 47124
rect 29204 47068 29214 47124
rect 30146 47068 30156 47124
rect 30212 47068 33684 47124
rect 44034 47068 44044 47124
rect 44100 47068 46956 47124
rect 47012 47068 48748 47124
rect 48804 47068 49756 47124
rect 49812 47068 49822 47124
rect 50978 47068 50988 47124
rect 51044 47068 51996 47124
rect 52052 47068 52668 47124
rect 52724 47068 52734 47124
rect 58146 47068 58156 47124
rect 58212 47068 60000 47124
rect 15092 47012 15148 47068
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 33628 47012 33684 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 59200 47040 60000 47068
rect 11676 46956 13020 47012
rect 13076 46956 13356 47012
rect 13412 46956 13422 47012
rect 13570 46956 13580 47012
rect 13636 46956 15148 47012
rect 16034 46956 16044 47012
rect 16100 46956 18172 47012
rect 18228 46956 18238 47012
rect 18722 46956 18732 47012
rect 18788 46956 19516 47012
rect 19572 46956 19582 47012
rect 21858 46956 21868 47012
rect 21924 46956 27244 47012
rect 27300 46956 27310 47012
rect 27458 46956 27468 47012
rect 27524 46956 28700 47012
rect 28756 46956 28766 47012
rect 29810 46956 29820 47012
rect 29876 46956 32172 47012
rect 32228 46956 32238 47012
rect 33618 46956 33628 47012
rect 33684 46956 33694 47012
rect 35522 46956 35532 47012
rect 35588 46956 36764 47012
rect 36820 46956 36830 47012
rect 38434 46956 38444 47012
rect 38500 46956 38780 47012
rect 38836 46956 41916 47012
rect 41972 46956 41982 47012
rect 44146 46956 44156 47012
rect 44212 46956 46060 47012
rect 46116 46956 46126 47012
rect 16268 46844 16492 46900
rect 16548 46844 16558 46900
rect 16818 46844 16828 46900
rect 16884 46844 18508 46900
rect 18564 46844 18574 46900
rect 19394 46844 19404 46900
rect 19460 46844 24220 46900
rect 24276 46844 27524 46900
rect 27682 46844 27692 46900
rect 27748 46844 28924 46900
rect 28980 46844 28990 46900
rect 29586 46844 29596 46900
rect 29652 46844 30044 46900
rect 30100 46844 30110 46900
rect 32946 46844 32956 46900
rect 33012 46844 33180 46900
rect 33236 46844 33246 46900
rect 40114 46844 40124 46900
rect 40180 46844 41580 46900
rect 41636 46844 41646 46900
rect 45154 46844 45164 46900
rect 45220 46844 45836 46900
rect 45892 46844 45902 46900
rect 16268 46788 16324 46844
rect 27468 46788 27524 46844
rect 14018 46732 14028 46788
rect 14084 46732 16268 46788
rect 16324 46732 16334 46788
rect 20514 46732 20524 46788
rect 20580 46732 21084 46788
rect 21140 46732 21150 46788
rect 23986 46732 23996 46788
rect 24052 46732 27132 46788
rect 27188 46732 27198 46788
rect 27458 46732 27468 46788
rect 27524 46732 30156 46788
rect 30212 46732 30222 46788
rect 49074 46732 49084 46788
rect 49140 46732 50316 46788
rect 50372 46732 50382 46788
rect 9202 46620 9212 46676
rect 9268 46620 9660 46676
rect 9716 46620 10332 46676
rect 10388 46620 10398 46676
rect 11974 46620 12012 46676
rect 12068 46620 12078 46676
rect 17042 46620 17052 46676
rect 17108 46620 17612 46676
rect 17668 46620 17678 46676
rect 18162 46620 18172 46676
rect 18228 46620 23772 46676
rect 23828 46620 23838 46676
rect 24882 46620 24892 46676
rect 24948 46620 26236 46676
rect 26292 46620 26302 46676
rect 26422 46620 26460 46676
rect 26516 46620 26526 46676
rect 26674 46620 26684 46676
rect 26740 46620 26778 46676
rect 27234 46620 27244 46676
rect 27300 46620 28476 46676
rect 28532 46620 28542 46676
rect 28690 46620 28700 46676
rect 28756 46620 29260 46676
rect 29316 46620 31388 46676
rect 31444 46620 31454 46676
rect 36194 46620 36204 46676
rect 36260 46620 39900 46676
rect 39956 46620 40908 46676
rect 40964 46620 40974 46676
rect 41234 46620 41244 46676
rect 41300 46620 42252 46676
rect 42308 46620 42924 46676
rect 42980 46620 42990 46676
rect 52322 46620 52332 46676
rect 52388 46620 53564 46676
rect 53620 46620 53630 46676
rect 6850 46508 6860 46564
rect 6916 46508 6972 46564
rect 7028 46508 7038 46564
rect 11890 46508 11900 46564
rect 11956 46508 12348 46564
rect 12404 46508 12414 46564
rect 15250 46508 15260 46564
rect 15316 46508 16492 46564
rect 16548 46508 23548 46564
rect 25554 46508 25564 46564
rect 25620 46508 26572 46564
rect 26628 46508 28588 46564
rect 28644 46508 33852 46564
rect 33908 46508 33918 46564
rect 36978 46508 36988 46564
rect 37044 46508 37996 46564
rect 38052 46508 38444 46564
rect 38500 46508 38510 46564
rect 23492 46452 23548 46508
rect 7634 46396 7644 46452
rect 7700 46396 8540 46452
rect 8596 46396 8606 46452
rect 8866 46396 8876 46452
rect 8932 46396 18732 46452
rect 18788 46396 20188 46452
rect 20244 46396 20254 46452
rect 23492 46396 26236 46452
rect 26292 46396 26796 46452
rect 26852 46396 26862 46452
rect 27010 46396 27020 46452
rect 27076 46396 27468 46452
rect 27524 46396 29596 46452
rect 29652 46396 29662 46452
rect 15922 46284 15932 46340
rect 15988 46284 23884 46340
rect 23940 46284 23950 46340
rect 24658 46284 24668 46340
rect 24724 46284 29260 46340
rect 29316 46284 29326 46340
rect 29474 46284 29484 46340
rect 29540 46284 29932 46340
rect 29988 46284 29998 46340
rect 30258 46284 30268 46340
rect 30324 46284 30828 46340
rect 30884 46284 30894 46340
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 16818 46172 16828 46228
rect 16884 46172 17836 46228
rect 17892 46172 17902 46228
rect 20290 46172 20300 46228
rect 20356 46172 21868 46228
rect 21924 46172 21934 46228
rect 25778 46172 25788 46228
rect 25844 46172 34076 46228
rect 34132 46172 34142 46228
rect 11554 46060 11564 46116
rect 11620 46060 18732 46116
rect 18788 46060 19740 46116
rect 19796 46060 19806 46116
rect 20402 46060 20412 46116
rect 20468 46060 21308 46116
rect 21364 46060 21374 46116
rect 22082 46060 22092 46116
rect 22148 46060 22764 46116
rect 22820 46060 22830 46116
rect 24770 46060 24780 46116
rect 24836 46060 25228 46116
rect 25284 46060 25294 46116
rect 28550 46060 28588 46116
rect 28644 46060 32284 46116
rect 32340 46060 32350 46116
rect 32834 46060 32844 46116
rect 32900 46060 41244 46116
rect 41300 46060 42140 46116
rect 42196 46060 42206 46116
rect 12898 45948 12908 46004
rect 12964 45948 15484 46004
rect 15540 45948 15550 46004
rect 18722 45948 18732 46004
rect 18788 45948 20860 46004
rect 20916 45948 20926 46004
rect 23846 45948 23884 46004
rect 23940 45948 23950 46004
rect 28018 45948 28028 46004
rect 28084 45948 28252 46004
rect 28308 45948 29372 46004
rect 29428 45948 29438 46004
rect 29922 45948 29932 46004
rect 29988 45948 30044 46004
rect 30100 45948 30110 46004
rect 48066 45948 48076 46004
rect 48132 45948 48748 46004
rect 48804 45948 48814 46004
rect 7186 45836 7196 45892
rect 7252 45836 8876 45892
rect 8932 45836 9884 45892
rect 9940 45836 10444 45892
rect 10500 45836 10510 45892
rect 11666 45836 11676 45892
rect 11732 45836 18956 45892
rect 19012 45836 22428 45892
rect 22484 45836 26572 45892
rect 26628 45836 26638 45892
rect 29474 45836 29484 45892
rect 29540 45836 31500 45892
rect 31556 45836 31566 45892
rect 34262 45836 34300 45892
rect 34356 45836 34366 45892
rect 6290 45724 6300 45780
rect 6356 45724 7644 45780
rect 7700 45724 7710 45780
rect 8754 45724 8764 45780
rect 8820 45724 11788 45780
rect 11844 45724 11854 45780
rect 14130 45724 14140 45780
rect 14196 45724 19236 45780
rect 19394 45724 19404 45780
rect 19460 45724 19740 45780
rect 19796 45724 21644 45780
rect 21700 45724 21710 45780
rect 23650 45724 23660 45780
rect 23716 45724 24444 45780
rect 24500 45724 24510 45780
rect 25666 45724 25676 45780
rect 25732 45724 27020 45780
rect 27076 45724 28700 45780
rect 28756 45724 28766 45780
rect 28914 45724 28924 45780
rect 28980 45724 29148 45780
rect 29204 45724 30380 45780
rect 30436 45724 30446 45780
rect 36642 45724 36652 45780
rect 36708 45724 39228 45780
rect 39284 45724 40012 45780
rect 40068 45724 40078 45780
rect 41906 45724 41916 45780
rect 41972 45724 48748 45780
rect 48804 45724 49196 45780
rect 49252 45724 49644 45780
rect 49700 45724 49710 45780
rect 19180 45668 19236 45724
rect 6066 45612 6076 45668
rect 6132 45612 6524 45668
rect 6580 45612 6590 45668
rect 9426 45612 9436 45668
rect 9492 45612 15148 45668
rect 19170 45612 19180 45668
rect 19236 45612 20076 45668
rect 20132 45612 20142 45668
rect 22754 45612 22764 45668
rect 22820 45612 23436 45668
rect 23492 45612 25340 45668
rect 25396 45612 25406 45668
rect 27346 45612 27356 45668
rect 27412 45612 32620 45668
rect 32676 45612 32686 45668
rect 38770 45612 38780 45668
rect 38836 45612 39788 45668
rect 39844 45612 39854 45668
rect 15092 45556 15148 45612
rect 8082 45500 8092 45556
rect 8148 45500 13804 45556
rect 13860 45500 13870 45556
rect 15092 45500 17388 45556
rect 17444 45500 17500 45556
rect 17556 45500 17566 45556
rect 20962 45500 20972 45556
rect 21028 45500 22204 45556
rect 22260 45500 22270 45556
rect 28802 45500 28812 45556
rect 28868 45500 29260 45556
rect 29316 45500 29326 45556
rect 31714 45500 31724 45556
rect 31780 45500 36876 45556
rect 36932 45500 36942 45556
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 9538 45388 9548 45444
rect 9604 45388 9614 45444
rect 14130 45388 14140 45444
rect 14196 45388 14812 45444
rect 14868 45388 14878 45444
rect 18050 45388 18060 45444
rect 18116 45388 19180 45444
rect 19236 45388 19246 45444
rect 21522 45388 21532 45444
rect 21588 45388 21924 45444
rect 23986 45388 23996 45444
rect 24052 45388 24668 45444
rect 24724 45388 25340 45444
rect 25396 45388 26572 45444
rect 26628 45388 26638 45444
rect 26898 45388 26908 45444
rect 26964 45388 27356 45444
rect 27412 45388 27422 45444
rect 27682 45388 27692 45444
rect 27748 45388 29932 45444
rect 29988 45388 29998 45444
rect 30482 45388 30492 45444
rect 30548 45388 32508 45444
rect 32564 45388 32574 45444
rect 39330 45388 39340 45444
rect 39396 45388 42476 45444
rect 42532 45388 42542 45444
rect 9548 45332 9604 45388
rect 21868 45332 21924 45388
rect 9548 45276 11228 45332
rect 11284 45276 11788 45332
rect 11844 45276 11854 45332
rect 19618 45276 19628 45332
rect 19684 45276 21532 45332
rect 21588 45276 21598 45332
rect 21868 45276 35364 45332
rect 48402 45276 48412 45332
rect 48468 45276 49308 45332
rect 49364 45276 49374 45332
rect 16706 45164 16716 45220
rect 16772 45164 18284 45220
rect 18340 45164 18350 45220
rect 19506 45164 19516 45220
rect 19572 45164 19740 45220
rect 19796 45164 19806 45220
rect 20178 45164 20188 45220
rect 20244 45164 22652 45220
rect 22708 45164 24444 45220
rect 24500 45164 24510 45220
rect 24770 45164 24780 45220
rect 24836 45164 25452 45220
rect 25508 45164 25518 45220
rect 28354 45164 28364 45220
rect 28420 45164 29708 45220
rect 29764 45164 29774 45220
rect 30146 45164 30156 45220
rect 30212 45164 33404 45220
rect 33460 45164 34076 45220
rect 34132 45164 34142 45220
rect 24444 45108 24500 45164
rect 35308 45108 35364 45276
rect 43362 45164 43372 45220
rect 43428 45164 45164 45220
rect 45220 45164 45230 45220
rect 45714 45164 45724 45220
rect 45780 45164 46844 45220
rect 46900 45164 46910 45220
rect 47730 45164 47740 45220
rect 47796 45164 48972 45220
rect 49028 45164 50316 45220
rect 50372 45164 50382 45220
rect 9986 45052 9996 45108
rect 10052 45052 13356 45108
rect 13412 45052 19964 45108
rect 20020 45052 20030 45108
rect 24444 45052 25116 45108
rect 25172 45052 25182 45108
rect 26236 45052 28476 45108
rect 28532 45052 28542 45108
rect 28802 45052 28812 45108
rect 28868 45052 31164 45108
rect 31220 45052 31230 45108
rect 32498 45052 32508 45108
rect 32564 45052 33852 45108
rect 33908 45052 33918 45108
rect 35298 45052 35308 45108
rect 35364 45052 35374 45108
rect 45378 45052 45388 45108
rect 45444 45052 47068 45108
rect 47124 45052 47134 45108
rect 47394 45052 47404 45108
rect 47460 45052 48748 45108
rect 48804 45052 48814 45108
rect 26236 44996 26292 45052
rect 46732 44996 46788 45052
rect 7858 44940 7868 44996
rect 7924 44940 13020 44996
rect 13076 44940 21196 44996
rect 21252 44940 21262 44996
rect 25890 44940 25900 44996
rect 25956 44940 26236 44996
rect 26292 44940 26302 44996
rect 28018 44940 28028 44996
rect 28084 44940 34524 44996
rect 34580 44940 34590 44996
rect 46722 44940 46732 44996
rect 46788 44940 46798 44996
rect 49970 44940 49980 44996
rect 50036 44940 50764 44996
rect 50820 44940 50830 44996
rect 13766 44828 13804 44884
rect 13860 44828 13870 44884
rect 15474 44828 15484 44884
rect 15540 44828 15708 44884
rect 15764 44828 16828 44884
rect 16884 44828 16894 44884
rect 19058 44828 19068 44884
rect 19124 44828 20524 44884
rect 20580 44828 27468 44884
rect 27524 44828 27534 44884
rect 28364 44828 34188 44884
rect 34244 44828 34748 44884
rect 34804 44828 34814 44884
rect 36418 44828 36428 44884
rect 36484 44828 43484 44884
rect 43540 44828 44940 44884
rect 44996 44828 45276 44884
rect 45332 44828 45342 44884
rect 46610 44828 46620 44884
rect 46676 44828 47180 44884
rect 47236 44828 47246 44884
rect 28364 44772 28420 44828
rect 19282 44716 19292 44772
rect 19348 44716 28420 44772
rect 28998 44716 29036 44772
rect 29092 44716 29102 44772
rect 33394 44716 33404 44772
rect 33460 44716 34300 44772
rect 34356 44716 34366 44772
rect 40114 44716 40124 44772
rect 40180 44716 41020 44772
rect 41076 44716 41086 44772
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 15810 44604 15820 44660
rect 15876 44604 17724 44660
rect 17780 44604 23884 44660
rect 23940 44604 25228 44660
rect 25284 44604 25294 44660
rect 14802 44492 14812 44548
rect 14868 44492 16716 44548
rect 16772 44492 16782 44548
rect 19506 44492 19516 44548
rect 19572 44492 23436 44548
rect 23492 44492 23502 44548
rect 24518 44492 24556 44548
rect 24612 44492 24622 44548
rect 28578 44492 28588 44548
rect 28644 44492 28700 44548
rect 28756 44492 29260 44548
rect 29316 44492 29326 44548
rect 31378 44492 31388 44548
rect 31444 44492 32284 44548
rect 32340 44492 32350 44548
rect 41346 44492 41356 44548
rect 41412 44492 47292 44548
rect 47348 44492 47516 44548
rect 47572 44492 47582 44548
rect 59200 44436 60000 44464
rect 11778 44380 11788 44436
rect 11844 44380 12684 44436
rect 12740 44380 12750 44436
rect 15474 44380 15484 44436
rect 15540 44380 18844 44436
rect 18900 44380 23772 44436
rect 23828 44380 23838 44436
rect 24882 44380 24892 44436
rect 24948 44380 27636 44436
rect 28690 44380 28700 44436
rect 28756 44380 29372 44436
rect 29428 44380 29438 44436
rect 31154 44380 31164 44436
rect 31220 44380 32732 44436
rect 32788 44380 33068 44436
rect 33124 44380 33134 44436
rect 34738 44380 34748 44436
rect 34804 44380 37100 44436
rect 37156 44380 37166 44436
rect 38210 44380 38220 44436
rect 38276 44380 50652 44436
rect 50708 44380 50988 44436
rect 51044 44380 51054 44436
rect 57922 44380 57932 44436
rect 57988 44380 60000 44436
rect 12898 44268 12908 44324
rect 12964 44268 14028 44324
rect 14084 44268 14094 44324
rect 15698 44268 15708 44324
rect 15764 44268 16380 44324
rect 16436 44268 18956 44324
rect 19012 44268 19516 44324
rect 19572 44268 19582 44324
rect 19842 44268 19852 44324
rect 19908 44268 21308 44324
rect 21364 44268 21374 44324
rect 21858 44268 21868 44324
rect 21924 44268 22988 44324
rect 23044 44268 24108 44324
rect 24164 44268 24174 44324
rect 24546 44268 24556 44324
rect 24612 44268 25004 44324
rect 25060 44268 25070 44324
rect 26450 44268 26460 44324
rect 26516 44268 26796 44324
rect 26852 44268 26862 44324
rect 13580 44156 16268 44212
rect 16324 44156 16334 44212
rect 16818 44156 16828 44212
rect 16884 44156 17276 44212
rect 17332 44156 17724 44212
rect 17780 44156 17790 44212
rect 19618 44156 19628 44212
rect 19684 44156 19964 44212
rect 20020 44156 20524 44212
rect 20580 44156 20590 44212
rect 23100 44156 26460 44212
rect 26516 44156 26908 44212
rect 13580 44100 13636 44156
rect 23100 44100 23156 44156
rect 7858 44044 7868 44100
rect 7924 44044 13580 44100
rect 13636 44044 13646 44100
rect 13794 44044 13804 44100
rect 13860 44044 14028 44100
rect 14084 44044 14094 44100
rect 14438 44044 14476 44100
rect 14532 44044 14542 44100
rect 14690 44044 14700 44100
rect 14756 44044 15148 44100
rect 15204 44044 15214 44100
rect 20738 44044 20748 44100
rect 20804 44044 21868 44100
rect 21924 44044 21934 44100
rect 23062 44044 23100 44100
rect 23156 44044 23166 44100
rect 23538 44044 23548 44100
rect 23604 44044 25340 44100
rect 25396 44044 26012 44100
rect 26068 44044 26078 44100
rect 14028 43988 14084 44044
rect 26852 43988 26908 44156
rect 27580 44100 27636 44380
rect 59200 44352 60000 44380
rect 29446 44268 29484 44324
rect 29540 44268 29550 44324
rect 29698 44268 29708 44324
rect 29764 44268 30604 44324
rect 30660 44268 30670 44324
rect 30930 44268 30940 44324
rect 30996 44268 31836 44324
rect 31892 44268 31902 44324
rect 35074 44268 35084 44324
rect 35140 44268 35868 44324
rect 35924 44268 35934 44324
rect 37986 44268 37996 44324
rect 38052 44268 38332 44324
rect 38388 44268 39004 44324
rect 39060 44268 42700 44324
rect 42756 44268 42766 44324
rect 45266 44268 45276 44324
rect 45332 44268 45836 44324
rect 45892 44268 45902 44324
rect 53106 44268 53116 44324
rect 53172 44268 54572 44324
rect 54628 44268 54638 44324
rect 27794 44156 27804 44212
rect 27860 44156 29820 44212
rect 29876 44156 29886 44212
rect 33058 44156 33068 44212
rect 33124 44156 36764 44212
rect 36820 44156 37548 44212
rect 37604 44156 37614 44212
rect 27010 44044 27020 44100
rect 27076 44044 27114 44100
rect 27580 44044 33404 44100
rect 33460 44044 33470 44100
rect 33618 44044 33628 44100
rect 33684 44044 35756 44100
rect 35812 44044 36316 44100
rect 36372 44044 36382 44100
rect 41458 44044 41468 44100
rect 41524 44044 42028 44100
rect 42084 44044 42094 44100
rect 43474 44044 43484 44100
rect 43540 44044 44828 44100
rect 44884 44044 44894 44100
rect 10322 43932 10332 43988
rect 10388 43932 11228 43988
rect 11284 43932 11900 43988
rect 11956 43932 11966 43988
rect 14028 43932 15484 43988
rect 15540 43932 15550 43988
rect 17602 43932 17612 43988
rect 17668 43932 18060 43988
rect 18116 43932 18126 43988
rect 26852 43932 31612 43988
rect 31668 43932 31678 43988
rect 34150 43932 34188 43988
rect 34244 43932 34254 43988
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 12786 43820 12796 43876
rect 12852 43820 18956 43876
rect 19012 43820 19022 43876
rect 29260 43764 29316 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 32274 43820 32284 43876
rect 32340 43820 34524 43876
rect 34580 43820 34860 43876
rect 34916 43820 34926 43876
rect 8082 43708 8092 43764
rect 8148 43708 14700 43764
rect 14756 43708 14766 43764
rect 17714 43708 17724 43764
rect 17780 43708 20636 43764
rect 20692 43708 20702 43764
rect 29250 43708 29260 43764
rect 29316 43708 29326 43764
rect 29922 43708 29932 43764
rect 29988 43708 30156 43764
rect 30212 43708 31052 43764
rect 31108 43708 31118 43764
rect 31378 43708 31388 43764
rect 31444 43708 32844 43764
rect 32900 43708 32910 43764
rect 33954 43708 33964 43764
rect 34020 43708 34972 43764
rect 35028 43708 35038 43764
rect 46050 43708 46060 43764
rect 46116 43708 46732 43764
rect 46788 43708 48412 43764
rect 48468 43708 48478 43764
rect 48636 43708 50092 43764
rect 50148 43708 50158 43764
rect 48636 43652 48692 43708
rect 14354 43596 14364 43652
rect 14420 43596 15148 43652
rect 19394 43596 19404 43652
rect 19460 43596 19740 43652
rect 19796 43596 19806 43652
rect 20402 43596 20412 43652
rect 20468 43596 21084 43652
rect 21140 43596 21150 43652
rect 22278 43596 22316 43652
rect 22372 43596 22382 43652
rect 22866 43596 22876 43652
rect 22932 43596 22942 43652
rect 23426 43596 23436 43652
rect 23492 43596 24332 43652
rect 24388 43596 24398 43652
rect 24882 43596 24892 43652
rect 24948 43596 25788 43652
rect 25844 43596 25854 43652
rect 26086 43596 26124 43652
rect 26180 43596 27020 43652
rect 27076 43596 27580 43652
rect 27636 43596 28588 43652
rect 28644 43596 28654 43652
rect 29138 43596 29148 43652
rect 29204 43596 30044 43652
rect 30100 43596 30604 43652
rect 30660 43596 30670 43652
rect 33394 43596 33404 43652
rect 33460 43596 34636 43652
rect 34692 43596 34702 43652
rect 37426 43596 37436 43652
rect 37492 43596 38668 43652
rect 38724 43596 38734 43652
rect 41580 43596 48692 43652
rect 51202 43596 51212 43652
rect 51268 43596 51772 43652
rect 51828 43596 52220 43652
rect 52276 43596 52286 43652
rect 53890 43596 53900 43652
rect 53956 43596 54460 43652
rect 54516 43596 54526 43652
rect 15092 43540 15148 43596
rect 22876 43540 22932 43596
rect 6626 43484 6636 43540
rect 6692 43484 8204 43540
rect 8260 43484 9548 43540
rect 9604 43484 9614 43540
rect 14130 43484 14140 43540
rect 14196 43484 14924 43540
rect 14980 43484 14990 43540
rect 15092 43484 15596 43540
rect 15652 43484 16212 43540
rect 18386 43484 18396 43540
rect 18452 43484 22932 43540
rect 23874 43484 23884 43540
rect 23940 43484 25340 43540
rect 25396 43484 25406 43540
rect 16156 43316 16212 43484
rect 26124 43428 26180 43596
rect 26786 43484 26796 43540
rect 26852 43484 29036 43540
rect 29092 43484 29596 43540
rect 29652 43484 30380 43540
rect 30436 43484 30446 43540
rect 30706 43484 30716 43540
rect 30772 43484 36428 43540
rect 36484 43484 37548 43540
rect 37604 43484 37772 43540
rect 37828 43484 37838 43540
rect 39666 43484 39676 43540
rect 39732 43484 40348 43540
rect 40404 43484 40908 43540
rect 40964 43484 40974 43540
rect 41580 43428 41636 43596
rect 41794 43484 41804 43540
rect 41860 43484 42588 43540
rect 42644 43484 42654 43540
rect 42914 43484 42924 43540
rect 42980 43484 44380 43540
rect 44436 43484 44446 43540
rect 47730 43484 47740 43540
rect 47796 43484 49084 43540
rect 49140 43484 49150 43540
rect 51650 43484 51660 43540
rect 51716 43484 52332 43540
rect 52388 43484 52398 43540
rect 52882 43484 52892 43540
rect 52948 43484 54796 43540
rect 54852 43484 54862 43540
rect 55458 43484 55468 43540
rect 55524 43484 56812 43540
rect 56868 43484 56878 43540
rect 16370 43372 16380 43428
rect 16436 43372 17388 43428
rect 17444 43372 19740 43428
rect 19796 43372 19806 43428
rect 21634 43372 21644 43428
rect 21700 43372 22316 43428
rect 22372 43372 22382 43428
rect 22754 43372 22764 43428
rect 22820 43372 23212 43428
rect 23268 43372 26180 43428
rect 26338 43372 26348 43428
rect 26404 43372 28700 43428
rect 28756 43372 28766 43428
rect 33730 43372 33740 43428
rect 33796 43372 34860 43428
rect 34916 43372 34926 43428
rect 38546 43372 38556 43428
rect 38612 43372 41636 43428
rect 43474 43372 43484 43428
rect 43540 43372 46172 43428
rect 46228 43372 46238 43428
rect 16156 43260 18228 43316
rect 20850 43260 20860 43316
rect 20916 43260 21420 43316
rect 21476 43260 21486 43316
rect 21746 43260 21756 43316
rect 21812 43260 26908 43316
rect 28578 43260 28588 43316
rect 28644 43260 39340 43316
rect 39396 43260 39406 43316
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 18172 43092 18228 43260
rect 26852 43204 26908 43260
rect 21970 43148 21980 43204
rect 22036 43148 23884 43204
rect 23940 43148 23950 43204
rect 24098 43148 24108 43204
rect 24164 43148 25900 43204
rect 25956 43148 25966 43204
rect 26852 43148 28924 43204
rect 28980 43148 28990 43204
rect 32050 43148 32060 43204
rect 32116 43148 33404 43204
rect 33460 43148 33470 43204
rect 45042 43148 45052 43204
rect 45108 43148 45500 43204
rect 45556 43148 45566 43204
rect 18172 43036 25564 43092
rect 25620 43036 25630 43092
rect 25900 42980 25956 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 59200 43092 60000 43120
rect 27458 43036 27468 43092
rect 27524 43036 27804 43092
rect 27860 43036 27870 43092
rect 29026 43036 29036 43092
rect 29092 43036 29708 43092
rect 29764 43036 29774 43092
rect 57922 43036 57932 43092
rect 57988 43036 60000 43092
rect 59200 43008 60000 43036
rect 12674 42924 12684 42980
rect 12740 42924 16268 42980
rect 16324 42924 18564 42980
rect 18722 42924 18732 42980
rect 18788 42924 20412 42980
rect 20468 42924 20478 42980
rect 21532 42924 25844 42980
rect 25900 42924 26908 42980
rect 27346 42924 27356 42980
rect 27412 42924 29428 42980
rect 29586 42924 29596 42980
rect 29652 42924 30044 42980
rect 30100 42924 30110 42980
rect 30818 42924 30828 42980
rect 30884 42924 32060 42980
rect 32116 42924 32126 42980
rect 33170 42924 33180 42980
rect 33236 42924 34300 42980
rect 34356 42924 34366 42980
rect 36306 42924 36316 42980
rect 36372 42924 45388 42980
rect 45444 42924 45454 42980
rect 45826 42924 45836 42980
rect 45892 42924 49420 42980
rect 49476 42924 49980 42980
rect 50036 42924 50046 42980
rect 18508 42868 18564 42924
rect 21532 42868 21588 42924
rect 25788 42868 25844 42924
rect 26852 42868 26908 42924
rect 29372 42868 29428 42924
rect 12562 42812 12572 42868
rect 12628 42812 18060 42868
rect 18116 42812 18284 42868
rect 18340 42812 18350 42868
rect 18508 42812 20860 42868
rect 20916 42812 21532 42868
rect 21588 42812 21598 42868
rect 25788 42812 26348 42868
rect 26404 42812 26414 42868
rect 26562 42812 26572 42868
rect 26628 42812 26638 42868
rect 26852 42812 27468 42868
rect 27524 42812 27534 42868
rect 29372 42812 37996 42868
rect 38052 42812 38062 42868
rect 49858 42812 49868 42868
rect 49924 42812 51212 42868
rect 51268 42812 51278 42868
rect 10658 42700 10668 42756
rect 10724 42700 11564 42756
rect 11620 42700 11630 42756
rect 15698 42700 15708 42756
rect 15764 42700 18732 42756
rect 18788 42700 18798 42756
rect 23538 42700 23548 42756
rect 23604 42700 23884 42756
rect 23940 42700 24444 42756
rect 24500 42700 24510 42756
rect 26572 42644 26628 42812
rect 26786 42700 26796 42756
rect 26852 42700 27356 42756
rect 27412 42700 27422 42756
rect 27570 42700 27580 42756
rect 27636 42700 28700 42756
rect 28756 42700 28766 42756
rect 30146 42700 30156 42756
rect 30212 42700 30380 42756
rect 30436 42700 30446 42756
rect 31826 42700 31836 42756
rect 31892 42700 32396 42756
rect 32452 42700 32462 42756
rect 45266 42700 45276 42756
rect 45332 42700 49420 42756
rect 49476 42700 50092 42756
rect 50148 42700 50158 42756
rect 51762 42700 51772 42756
rect 51828 42700 53004 42756
rect 53060 42700 53070 42756
rect 8306 42588 8316 42644
rect 8372 42588 16156 42644
rect 16212 42588 16222 42644
rect 17042 42588 17052 42644
rect 17108 42588 19404 42644
rect 19460 42588 19470 42644
rect 19628 42588 22092 42644
rect 22148 42588 22158 42644
rect 26572 42588 31276 42644
rect 31332 42588 32508 42644
rect 32564 42588 32574 42644
rect 32722 42588 32732 42644
rect 32788 42588 35532 42644
rect 35588 42588 35598 42644
rect 36642 42588 36652 42644
rect 36708 42588 37884 42644
rect 37940 42588 37950 42644
rect 41906 42588 41916 42644
rect 41972 42588 42588 42644
rect 42644 42588 42924 42644
rect 42980 42588 43596 42644
rect 43652 42588 43662 42644
rect 0 42420 800 42448
rect 19628 42420 19684 42588
rect 21522 42476 21532 42532
rect 21588 42476 28252 42532
rect 28308 42476 28318 42532
rect 30706 42476 30716 42532
rect 30772 42476 31164 42532
rect 31220 42476 31612 42532
rect 31668 42476 31678 42532
rect 38546 42476 38556 42532
rect 38612 42476 38892 42532
rect 38948 42476 38958 42532
rect 48850 42476 48860 42532
rect 48916 42476 51548 42532
rect 51604 42476 51614 42532
rect 0 42364 1708 42420
rect 1764 42364 1774 42420
rect 17154 42364 17164 42420
rect 17220 42364 19684 42420
rect 24098 42364 24108 42420
rect 24164 42364 26796 42420
rect 26852 42364 26862 42420
rect 27906 42364 27916 42420
rect 27972 42364 30604 42420
rect 30660 42364 30670 42420
rect 46470 42364 46508 42420
rect 46564 42364 46574 42420
rect 0 42336 800 42364
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 11666 42252 11676 42308
rect 11732 42252 15260 42308
rect 15316 42252 15326 42308
rect 26338 42252 26348 42308
rect 26404 42252 26908 42308
rect 26964 42252 26974 42308
rect 35634 42252 35644 42308
rect 35700 42252 36652 42308
rect 36708 42252 36718 42308
rect 8530 42140 8540 42196
rect 8596 42140 11452 42196
rect 11508 42140 11518 42196
rect 14914 42140 14924 42196
rect 14980 42140 21756 42196
rect 21812 42140 21822 42196
rect 22194 42140 22204 42196
rect 22260 42140 24332 42196
rect 24388 42140 24398 42196
rect 26674 42140 26684 42196
rect 26740 42140 26796 42196
rect 26852 42140 26862 42196
rect 33730 42140 33740 42196
rect 33796 42140 34972 42196
rect 35028 42140 35038 42196
rect 48178 42140 48188 42196
rect 48244 42140 49084 42196
rect 49140 42140 49150 42196
rect 51874 42140 51884 42196
rect 51940 42140 52556 42196
rect 52612 42140 53452 42196
rect 53508 42140 53518 42196
rect 18946 42028 18956 42084
rect 19012 42028 19292 42084
rect 19348 42028 19964 42084
rect 20020 42028 21308 42084
rect 21364 42028 21374 42084
rect 22204 42028 22316 42084
rect 22372 42028 22382 42084
rect 23622 42028 23660 42084
rect 23716 42028 23726 42084
rect 25554 42028 25564 42084
rect 25620 42028 25900 42084
rect 25956 42028 28924 42084
rect 28980 42028 28990 42084
rect 31154 42028 31164 42084
rect 31220 42028 34860 42084
rect 34916 42028 34926 42084
rect 47506 42028 47516 42084
rect 47572 42028 48412 42084
rect 48468 42028 49308 42084
rect 49364 42028 49374 42084
rect 22204 41972 22260 42028
rect 23660 41972 23716 42028
rect 10322 41916 10332 41972
rect 10388 41916 10668 41972
rect 10724 41916 10734 41972
rect 11330 41916 11340 41972
rect 11396 41916 12124 41972
rect 12180 41916 12190 41972
rect 12450 41916 12460 41972
rect 12516 41916 13804 41972
rect 13860 41916 13870 41972
rect 14550 41916 14588 41972
rect 14644 41916 14654 41972
rect 14914 41916 14924 41972
rect 14980 41916 15148 41972
rect 17350 41916 17388 41972
rect 17444 41916 17454 41972
rect 19394 41916 19404 41972
rect 19460 41916 19740 41972
rect 19796 41916 22260 41972
rect 22418 41916 22428 41972
rect 22484 41916 23716 41972
rect 26852 41916 27356 41972
rect 27412 41916 27422 41972
rect 28354 41916 28364 41972
rect 28420 41916 29372 41972
rect 29428 41916 29438 41972
rect 29586 41916 29596 41972
rect 29652 41916 29820 41972
rect 29876 41916 30604 41972
rect 30660 41916 30670 41972
rect 30818 41916 30828 41972
rect 30884 41916 31500 41972
rect 31556 41916 31566 41972
rect 34178 41916 34188 41972
rect 34244 41916 35196 41972
rect 35252 41916 35262 41972
rect 40226 41916 40236 41972
rect 40292 41916 42028 41972
rect 42084 41916 42476 41972
rect 42532 41916 42542 41972
rect 45714 41916 45724 41972
rect 45780 41916 47292 41972
rect 47348 41916 47358 41972
rect 47842 41916 47852 41972
rect 47908 41916 48972 41972
rect 49028 41916 49038 41972
rect 49186 41916 49196 41972
rect 49252 41916 51212 41972
rect 51268 41916 51278 41972
rect 51426 41916 51436 41972
rect 51492 41916 52444 41972
rect 52500 41916 52510 41972
rect 12674 41804 12684 41860
rect 12740 41804 13356 41860
rect 13412 41804 13422 41860
rect 15092 41804 15148 41916
rect 15204 41804 15214 41860
rect 17490 41804 17500 41860
rect 17556 41804 18396 41860
rect 18452 41804 18462 41860
rect 22204 41748 22260 41916
rect 26852 41860 26908 41916
rect 28364 41860 28420 41916
rect 25666 41804 25676 41860
rect 25732 41804 26908 41860
rect 27010 41804 27020 41860
rect 27076 41804 28420 41860
rect 34962 41804 34972 41860
rect 35028 41804 37996 41860
rect 38052 41804 38062 41860
rect 7298 41692 7308 41748
rect 7364 41692 8204 41748
rect 8260 41692 8270 41748
rect 11106 41692 11116 41748
rect 11172 41692 22148 41748
rect 22204 41692 22652 41748
rect 22708 41692 22718 41748
rect 26562 41692 26572 41748
rect 26628 41692 28476 41748
rect 28532 41692 28542 41748
rect 46162 41692 46172 41748
rect 46228 41692 47292 41748
rect 47348 41692 47358 41748
rect 22092 41636 22148 41692
rect 17826 41580 17836 41636
rect 17892 41580 20188 41636
rect 20244 41580 21084 41636
rect 21140 41580 21150 41636
rect 22082 41580 22092 41636
rect 22148 41580 22158 41636
rect 22652 41580 24220 41636
rect 24276 41580 26460 41636
rect 26516 41580 26526 41636
rect 46498 41580 46508 41636
rect 46564 41580 46732 41636
rect 46788 41580 46798 41636
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 22652 41524 22708 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 16258 41468 16268 41524
rect 16324 41468 22708 41524
rect 22866 41468 22876 41524
rect 22932 41468 23436 41524
rect 23492 41468 34412 41524
rect 34468 41468 34478 41524
rect 17378 41356 17388 41412
rect 17444 41356 17948 41412
rect 18004 41356 18014 41412
rect 19282 41356 19292 41412
rect 19348 41356 19628 41412
rect 19684 41356 19694 41412
rect 22306 41356 22316 41412
rect 22372 41356 23100 41412
rect 23156 41356 26012 41412
rect 26068 41356 26078 41412
rect 26338 41356 26348 41412
rect 26404 41356 27804 41412
rect 27860 41356 27870 41412
rect 30034 41356 30044 41412
rect 30100 41356 31276 41412
rect 31332 41356 33628 41412
rect 33684 41356 33694 41412
rect 42018 41356 42028 41412
rect 42084 41356 47068 41412
rect 47124 41356 47134 41412
rect 1698 41244 1708 41300
rect 1764 41244 1774 41300
rect 15092 41244 15372 41300
rect 15428 41244 18284 41300
rect 18340 41244 18956 41300
rect 19012 41244 19022 41300
rect 21746 41244 21756 41300
rect 21812 41244 22540 41300
rect 22596 41244 22606 41300
rect 22764 41244 31388 41300
rect 31444 41244 31454 41300
rect 46610 41244 46620 41300
rect 46676 41244 48076 41300
rect 48132 41244 48142 41300
rect 49074 41244 49084 41300
rect 49140 41244 49980 41300
rect 50036 41244 50046 41300
rect 0 41076 800 41104
rect 1708 41076 1764 41244
rect 15092 41188 15148 41244
rect 22764 41188 22820 41244
rect 6626 41132 6636 41188
rect 6692 41132 7084 41188
rect 7140 41132 7150 41188
rect 9762 41132 9772 41188
rect 9828 41132 14364 41188
rect 14420 41132 15148 41188
rect 16258 41132 16268 41188
rect 16324 41132 17388 41188
rect 17444 41132 17454 41188
rect 18386 41132 18396 41188
rect 18452 41132 22820 41188
rect 25218 41132 25228 41188
rect 25284 41132 28588 41188
rect 28644 41132 28654 41188
rect 28812 41132 29708 41188
rect 29764 41132 31500 41188
rect 31556 41132 31566 41188
rect 39666 41132 39676 41188
rect 39732 41132 41692 41188
rect 41748 41132 41758 41188
rect 47618 41132 47628 41188
rect 47684 41132 48636 41188
rect 48692 41132 48702 41188
rect 28812 41076 28868 41132
rect 0 41020 1764 41076
rect 11330 41020 11340 41076
rect 11396 41020 12684 41076
rect 12740 41020 12750 41076
rect 17266 41020 17276 41076
rect 17332 41020 17724 41076
rect 17780 41020 17790 41076
rect 18732 41020 19292 41076
rect 19348 41020 19358 41076
rect 19618 41020 19628 41076
rect 19684 41020 20524 41076
rect 20580 41020 20590 41076
rect 20738 41020 20748 41076
rect 20804 41020 21196 41076
rect 21252 41020 22092 41076
rect 22148 41020 22158 41076
rect 24182 41020 24220 41076
rect 24276 41020 24286 41076
rect 24780 41020 25564 41076
rect 25620 41020 25630 41076
rect 28690 41020 28700 41076
rect 28756 41020 28868 41076
rect 34066 41020 34076 41076
rect 34132 41020 34748 41076
rect 34804 41020 34814 41076
rect 38658 41020 38668 41076
rect 38724 41020 47852 41076
rect 47908 41020 48748 41076
rect 48804 41020 48814 41076
rect 51762 41020 51772 41076
rect 51828 41020 53004 41076
rect 53060 41020 53070 41076
rect 54338 41020 54348 41076
rect 54404 41020 55132 41076
rect 55188 41020 55198 41076
rect 0 40992 800 41020
rect 18732 40964 18788 41020
rect 24780 40964 24836 41020
rect 9762 40908 9772 40964
rect 9828 40908 10556 40964
rect 10612 40908 11004 40964
rect 11060 40908 11070 40964
rect 11228 40908 18788 40964
rect 18844 40908 20076 40964
rect 20132 40908 20142 40964
rect 23426 40908 23436 40964
rect 23492 40908 24780 40964
rect 24836 40908 24846 40964
rect 25638 40908 25676 40964
rect 25732 40908 25742 40964
rect 26114 40908 26124 40964
rect 26180 40908 29036 40964
rect 29092 40908 29102 40964
rect 36530 40908 36540 40964
rect 36596 40908 37212 40964
rect 37268 40908 37278 40964
rect 46274 40908 46284 40964
rect 46340 40908 46732 40964
rect 46788 40908 46798 40964
rect 48178 40908 48188 40964
rect 48244 40908 50988 40964
rect 51044 40908 51054 40964
rect 11228 40852 11284 40908
rect 18844 40852 18900 40908
rect 6850 40796 6860 40852
rect 6916 40796 7420 40852
rect 7476 40796 7980 40852
rect 8036 40796 8046 40852
rect 9650 40796 9660 40852
rect 9716 40796 11284 40852
rect 13346 40796 13356 40852
rect 13412 40796 18844 40852
rect 18900 40796 18910 40852
rect 20738 40796 20748 40852
rect 20804 40796 21644 40852
rect 21700 40796 25340 40852
rect 25396 40796 25406 40852
rect 32162 40796 32172 40852
rect 32228 40796 32238 40852
rect 13356 40740 13412 40796
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 32172 40740 32228 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 8866 40684 8876 40740
rect 8932 40684 13412 40740
rect 16930 40684 16940 40740
rect 16996 40684 17276 40740
rect 17332 40684 17342 40740
rect 26852 40684 32228 40740
rect 26852 40628 26908 40684
rect 9874 40572 9884 40628
rect 9940 40572 12012 40628
rect 12068 40572 12078 40628
rect 14914 40572 14924 40628
rect 14980 40572 15148 40628
rect 15204 40572 16492 40628
rect 16548 40572 16558 40628
rect 19730 40572 19740 40628
rect 19796 40572 20748 40628
rect 20804 40572 20814 40628
rect 22166 40572 22204 40628
rect 22260 40572 22270 40628
rect 26562 40572 26572 40628
rect 26628 40572 26908 40628
rect 27356 40572 27916 40628
rect 27972 40572 27982 40628
rect 28354 40572 28364 40628
rect 28420 40572 29708 40628
rect 29764 40572 29774 40628
rect 30818 40572 30828 40628
rect 30884 40572 33068 40628
rect 33124 40572 36988 40628
rect 37044 40572 37054 40628
rect 41794 40572 41804 40628
rect 41860 40572 45612 40628
rect 45668 40572 45678 40628
rect 53666 40572 53676 40628
rect 53732 40572 54460 40628
rect 54516 40572 54526 40628
rect 7522 40460 7532 40516
rect 7588 40460 7598 40516
rect 10210 40460 10220 40516
rect 10276 40460 10892 40516
rect 10948 40460 10958 40516
rect 17714 40460 17724 40516
rect 17780 40460 21196 40516
rect 21252 40460 21262 40516
rect 22642 40460 22652 40516
rect 22708 40460 27132 40516
rect 27188 40460 27198 40516
rect 7532 40292 7588 40460
rect 10098 40348 10108 40404
rect 10164 40348 11452 40404
rect 11508 40348 11676 40404
rect 11732 40348 11742 40404
rect 14130 40348 14140 40404
rect 14196 40348 14700 40404
rect 14756 40348 16268 40404
rect 16324 40348 16334 40404
rect 19142 40348 19180 40404
rect 19236 40348 19246 40404
rect 24322 40348 24332 40404
rect 24388 40348 25788 40404
rect 25844 40348 25854 40404
rect 27356 40292 27412 40572
rect 28578 40460 28588 40516
rect 28644 40460 29596 40516
rect 29652 40460 29662 40516
rect 49410 40460 49420 40516
rect 49476 40460 50540 40516
rect 50596 40460 51660 40516
rect 51716 40460 51726 40516
rect 59200 40404 60000 40432
rect 31490 40348 31500 40404
rect 31556 40348 31948 40404
rect 32004 40348 32014 40404
rect 35074 40348 35084 40404
rect 35140 40348 38780 40404
rect 38836 40348 38846 40404
rect 46274 40348 46284 40404
rect 46340 40348 47068 40404
rect 55234 40348 55244 40404
rect 55300 40348 56924 40404
rect 56980 40348 56990 40404
rect 57922 40348 57932 40404
rect 57988 40348 60000 40404
rect 47012 40292 47068 40348
rect 59200 40320 60000 40348
rect 7532 40236 8988 40292
rect 9044 40236 10668 40292
rect 10724 40236 10734 40292
rect 12786 40236 12796 40292
rect 12852 40236 15820 40292
rect 15876 40236 15886 40292
rect 16930 40236 16940 40292
rect 16996 40236 17836 40292
rect 17892 40236 17902 40292
rect 18946 40236 18956 40292
rect 19012 40236 21308 40292
rect 21364 40236 21374 40292
rect 24658 40236 24668 40292
rect 24724 40236 25564 40292
rect 25620 40236 25630 40292
rect 27234 40236 27244 40292
rect 27300 40236 27412 40292
rect 27682 40236 27692 40292
rect 27748 40236 29148 40292
rect 29204 40236 29820 40292
rect 29876 40236 29886 40292
rect 30146 40236 30156 40292
rect 30212 40236 30222 40292
rect 47012 40236 47292 40292
rect 47348 40236 47358 40292
rect 55010 40236 55020 40292
rect 55076 40236 56812 40292
rect 56868 40236 56878 40292
rect 30156 40180 30212 40236
rect 8082 40124 8092 40180
rect 8148 40124 9212 40180
rect 9268 40124 9278 40180
rect 14802 40124 14812 40180
rect 14868 40124 17388 40180
rect 17444 40124 17454 40180
rect 24994 40124 25004 40180
rect 25060 40124 30212 40180
rect 31714 40124 31724 40180
rect 31780 40124 32060 40180
rect 32116 40124 32126 40180
rect 7298 40012 7308 40068
rect 7364 40012 8428 40068
rect 8484 40012 8494 40068
rect 14354 40012 14364 40068
rect 14420 40012 14700 40068
rect 14756 40012 20748 40068
rect 20804 40012 21644 40068
rect 21700 40012 21710 40068
rect 22418 40012 22428 40068
rect 22484 40012 23324 40068
rect 23380 40012 23390 40068
rect 33814 40012 33852 40068
rect 33908 40012 33918 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 14914 39900 14924 39956
rect 14980 39900 18956 39956
rect 19012 39900 19022 39956
rect 50754 39900 50764 39956
rect 50820 39900 51100 39956
rect 51156 39900 51166 39956
rect 20626 39788 20636 39844
rect 20692 39788 22652 39844
rect 22708 39788 22718 39844
rect 26002 39788 26012 39844
rect 26068 39788 27580 39844
rect 27636 39788 29484 39844
rect 29540 39788 29550 39844
rect 49074 39788 49084 39844
rect 49140 39788 49532 39844
rect 49588 39788 49598 39844
rect 20636 39732 20692 39788
rect 10658 39676 10668 39732
rect 10724 39676 13468 39732
rect 13524 39676 13534 39732
rect 14914 39676 14924 39732
rect 14980 39676 16268 39732
rect 16324 39676 16334 39732
rect 18386 39676 18396 39732
rect 18452 39676 20692 39732
rect 22418 39676 22428 39732
rect 22484 39676 23100 39732
rect 23156 39676 23166 39732
rect 23874 39676 23884 39732
rect 23940 39676 27692 39732
rect 27748 39676 27758 39732
rect 28018 39676 28028 39732
rect 28084 39676 32284 39732
rect 32340 39676 32350 39732
rect 33506 39676 33516 39732
rect 33572 39676 36092 39732
rect 36148 39676 36158 39732
rect 27692 39620 27748 39676
rect 6626 39564 6636 39620
rect 6692 39564 7308 39620
rect 7364 39564 7374 39620
rect 8194 39564 8204 39620
rect 8260 39564 9996 39620
rect 10052 39564 11900 39620
rect 11956 39564 11966 39620
rect 15810 39564 15820 39620
rect 15876 39564 16604 39620
rect 16660 39564 16670 39620
rect 17938 39564 17948 39620
rect 18004 39564 19292 39620
rect 19348 39564 19358 39620
rect 22082 39564 22092 39620
rect 22148 39564 25452 39620
rect 25508 39564 25518 39620
rect 27692 39564 29148 39620
rect 29204 39564 29214 39620
rect 29922 39564 29932 39620
rect 29988 39564 31948 39620
rect 32004 39564 32014 39620
rect 34402 39564 34412 39620
rect 34468 39564 34860 39620
rect 34916 39564 34926 39620
rect 46050 39564 46060 39620
rect 46116 39564 48412 39620
rect 48468 39564 49756 39620
rect 49812 39564 49822 39620
rect 14018 39452 14028 39508
rect 14084 39452 14812 39508
rect 14868 39452 16940 39508
rect 16996 39452 17006 39508
rect 17826 39452 17836 39508
rect 17892 39452 19740 39508
rect 19796 39452 19806 39508
rect 20188 39452 25116 39508
rect 25172 39452 25340 39508
rect 25396 39452 25406 39508
rect 25666 39452 25676 39508
rect 25732 39452 35756 39508
rect 35812 39452 35822 39508
rect 48962 39452 48972 39508
rect 49028 39452 49644 39508
rect 49700 39452 50092 39508
rect 50148 39452 50158 39508
rect 50978 39452 50988 39508
rect 51044 39452 53228 39508
rect 53284 39452 53294 39508
rect 16940 39396 16996 39452
rect 7522 39340 7532 39396
rect 7588 39340 8092 39396
rect 8148 39340 8158 39396
rect 11554 39340 11564 39396
rect 11620 39340 16884 39396
rect 16940 39340 18284 39396
rect 18340 39340 18350 39396
rect 18918 39340 18956 39396
rect 19012 39340 19022 39396
rect 16828 39284 16884 39340
rect 7970 39228 7980 39284
rect 8036 39228 8428 39284
rect 8484 39228 8494 39284
rect 14662 39228 14700 39284
rect 14756 39228 14766 39284
rect 16828 39228 19180 39284
rect 19236 39228 19516 39284
rect 19572 39228 19582 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 7858 39116 7868 39172
rect 7924 39116 10332 39172
rect 10388 39116 14924 39172
rect 14980 39116 14990 39172
rect 0 39060 800 39088
rect 20188 39060 20244 39452
rect 22194 39340 22204 39396
rect 22260 39340 22652 39396
rect 22708 39340 22718 39396
rect 23874 39340 23884 39396
rect 23940 39340 23996 39396
rect 24052 39340 24062 39396
rect 26898 39340 26908 39396
rect 26964 39340 28028 39396
rect 28084 39340 28094 39396
rect 28578 39340 28588 39396
rect 28644 39340 29260 39396
rect 29316 39340 29326 39396
rect 34290 39340 34300 39396
rect 34356 39340 35980 39396
rect 36036 39340 36046 39396
rect 39890 39340 39900 39396
rect 39956 39340 41804 39396
rect 41860 39340 41870 39396
rect 42690 39340 42700 39396
rect 42756 39340 46284 39396
rect 46340 39340 46620 39396
rect 46676 39340 46686 39396
rect 46834 39340 46844 39396
rect 46900 39340 48636 39396
rect 48692 39340 49868 39396
rect 49924 39340 49934 39396
rect 20738 39228 20748 39284
rect 20804 39228 23324 39284
rect 23380 39228 31724 39284
rect 31780 39228 31790 39284
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 24210 39116 24220 39172
rect 24276 39116 32060 39172
rect 32116 39116 33516 39172
rect 33572 39116 33852 39172
rect 33908 39116 33918 39172
rect 41570 39116 41580 39172
rect 41636 39116 42364 39172
rect 42420 39116 43036 39172
rect 43092 39116 43102 39172
rect 0 39004 1708 39060
rect 1764 39004 1774 39060
rect 11890 39004 11900 39060
rect 11956 39004 12572 39060
rect 12628 39004 12638 39060
rect 15250 39004 15260 39060
rect 15316 39004 20244 39060
rect 21074 39004 21084 39060
rect 21140 39004 24108 39060
rect 24164 39004 25676 39060
rect 25732 39004 25742 39060
rect 26002 39004 26012 39060
rect 26068 39004 26796 39060
rect 26852 39004 26862 39060
rect 33394 39004 33404 39060
rect 33460 39004 33628 39060
rect 33684 39004 36316 39060
rect 36372 39004 36382 39060
rect 43586 39004 43596 39060
rect 43652 39004 45948 39060
rect 46004 39004 46014 39060
rect 47842 39004 47852 39060
rect 47908 39004 48972 39060
rect 49028 39004 49308 39060
rect 49364 39004 49374 39060
rect 49634 39004 49644 39060
rect 49700 39004 51100 39060
rect 51156 39004 51166 39060
rect 53218 39004 53228 39060
rect 53284 39004 54124 39060
rect 54180 39004 54572 39060
rect 54628 39004 54638 39060
rect 0 38976 800 39004
rect 15260 38948 15316 39004
rect 9986 38892 9996 38948
rect 10052 38892 14364 38948
rect 14420 38892 14430 38948
rect 15036 38892 15316 38948
rect 16940 38892 20860 38948
rect 20916 38892 23772 38948
rect 23828 38892 23838 38948
rect 34850 38892 34860 38948
rect 34916 38892 35756 38948
rect 35812 38892 35822 38948
rect 42578 38892 42588 38948
rect 42644 38892 45612 38948
rect 45668 38892 45678 38948
rect 50082 38892 50092 38948
rect 50148 38892 50540 38948
rect 50596 38892 50606 38948
rect 15036 38836 15092 38892
rect 12226 38780 12236 38836
rect 12292 38780 15092 38836
rect 16940 38724 16996 38892
rect 17154 38780 17164 38836
rect 17220 38780 17948 38836
rect 18004 38780 18014 38836
rect 22306 38780 22316 38836
rect 22372 38780 26124 38836
rect 26180 38780 26190 38836
rect 27458 38780 27468 38836
rect 27524 38780 29484 38836
rect 29540 38780 34188 38836
rect 34244 38780 34254 38836
rect 41570 38780 41580 38836
rect 41636 38780 42140 38836
rect 42196 38780 43260 38836
rect 43316 38780 43326 38836
rect 45154 38780 45164 38836
rect 45220 38780 46396 38836
rect 46452 38780 46462 38836
rect 51874 38780 51884 38836
rect 51940 38780 53116 38836
rect 53172 38780 54012 38836
rect 54068 38780 54078 38836
rect 11218 38668 11228 38724
rect 11284 38668 11788 38724
rect 11844 38668 11854 38724
rect 13122 38668 13132 38724
rect 13188 38668 14588 38724
rect 14644 38668 16996 38724
rect 19506 38668 19516 38724
rect 19572 38668 19964 38724
rect 20020 38668 23100 38724
rect 23156 38668 23166 38724
rect 23436 38668 23884 38724
rect 23940 38668 23950 38724
rect 32050 38668 32060 38724
rect 32116 38668 32508 38724
rect 32564 38668 34412 38724
rect 34468 38668 34478 38724
rect 35634 38668 35644 38724
rect 35700 38668 38332 38724
rect 38388 38668 38398 38724
rect 39218 38668 39228 38724
rect 39284 38668 48748 38724
rect 48804 38668 48814 38724
rect 23436 38612 23492 38668
rect 15362 38556 15372 38612
rect 15428 38556 15438 38612
rect 19058 38556 19068 38612
rect 19124 38556 19236 38612
rect 20290 38556 20300 38612
rect 20356 38556 20636 38612
rect 20692 38556 20702 38612
rect 22194 38556 22204 38612
rect 22260 38556 23492 38612
rect 23762 38556 23772 38612
rect 23828 38556 24892 38612
rect 24948 38556 24958 38612
rect 29222 38556 29260 38612
rect 29316 38556 29326 38612
rect 15372 38500 15428 38556
rect 19180 38500 19236 38556
rect 15372 38444 17500 38500
rect 17556 38444 17566 38500
rect 19170 38444 19180 38500
rect 19236 38444 19246 38500
rect 21522 38444 21532 38500
rect 21588 38444 26908 38500
rect 29026 38444 29036 38500
rect 29092 38444 32844 38500
rect 32900 38444 32910 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 26852 38388 26908 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 14242 38332 14252 38388
rect 14308 38332 25228 38388
rect 25284 38332 25294 38388
rect 26852 38332 30940 38388
rect 30996 38332 31006 38388
rect 11778 38220 11788 38276
rect 11844 38220 25900 38276
rect 25956 38220 25966 38276
rect 26226 38220 26236 38276
rect 26292 38220 30548 38276
rect 33282 38220 33292 38276
rect 33348 38220 41580 38276
rect 41636 38220 41646 38276
rect 30492 38164 30548 38220
rect 16146 38108 16156 38164
rect 16212 38108 17164 38164
rect 17220 38108 17230 38164
rect 19282 38108 19292 38164
rect 19348 38108 21084 38164
rect 21140 38108 21150 38164
rect 22278 38108 22316 38164
rect 22372 38108 22382 38164
rect 26852 38108 27692 38164
rect 27748 38108 27758 38164
rect 28130 38108 28140 38164
rect 28196 38108 30156 38164
rect 30212 38108 30222 38164
rect 30492 38108 34188 38164
rect 34244 38108 34254 38164
rect 26852 38052 26908 38108
rect 30156 38052 30212 38108
rect 16258 37996 16268 38052
rect 16324 37996 17836 38052
rect 17892 37996 17902 38052
rect 18722 37996 18732 38052
rect 18788 37996 19628 38052
rect 19684 37996 19694 38052
rect 20738 37996 20748 38052
rect 20804 37996 22876 38052
rect 22932 37996 23436 38052
rect 23492 37996 23502 38052
rect 26562 37996 26572 38052
rect 26628 37996 26908 38052
rect 28578 37996 28588 38052
rect 28644 37996 29260 38052
rect 29316 37996 29326 38052
rect 29474 37996 29484 38052
rect 29540 37996 29578 38052
rect 30156 37996 31164 38052
rect 31220 37996 31230 38052
rect 33030 37996 33068 38052
rect 33124 37996 33134 38052
rect 42802 37996 42812 38052
rect 42868 37996 43260 38052
rect 43316 37996 43326 38052
rect 53442 37996 53452 38052
rect 53508 37996 54796 38052
rect 54852 37996 54862 38052
rect 8306 37884 8316 37940
rect 8372 37884 10220 37940
rect 10276 37884 10286 37940
rect 18498 37884 18508 37940
rect 18564 37884 19628 37940
rect 19684 37884 19694 37940
rect 22082 37884 22092 37940
rect 22148 37884 22988 37940
rect 23044 37884 23054 37940
rect 26012 37884 27132 37940
rect 27188 37884 27198 37940
rect 28242 37884 28252 37940
rect 28308 37884 29708 37940
rect 29764 37884 29774 37940
rect 29932 37884 36092 37940
rect 36148 37884 37548 37940
rect 37604 37884 37614 37940
rect 41346 37884 41356 37940
rect 41412 37884 42252 37940
rect 42308 37884 42318 37940
rect 26012 37828 26068 37884
rect 10546 37772 10556 37828
rect 10612 37772 13468 37828
rect 13524 37772 15484 37828
rect 15540 37772 15550 37828
rect 17938 37772 17948 37828
rect 18004 37772 20188 37828
rect 20244 37772 21308 37828
rect 21364 37772 21374 37828
rect 23538 37772 23548 37828
rect 23604 37772 24220 37828
rect 24276 37772 26012 37828
rect 26068 37772 26078 37828
rect 26898 37772 26908 37828
rect 26964 37772 28028 37828
rect 28084 37772 28924 37828
rect 28980 37772 28990 37828
rect 29932 37716 29988 37884
rect 34290 37772 34300 37828
rect 34356 37772 35756 37828
rect 35812 37772 35822 37828
rect 37874 37772 37884 37828
rect 37940 37772 39004 37828
rect 39060 37772 39070 37828
rect 59200 37716 60000 37744
rect 21858 37660 21868 37716
rect 21924 37660 26796 37716
rect 26852 37660 27020 37716
rect 27076 37660 27086 37716
rect 27682 37660 27692 37716
rect 27748 37660 29988 37716
rect 30146 37660 30156 37716
rect 30212 37660 32620 37716
rect 32676 37660 32686 37716
rect 35970 37660 35980 37716
rect 36036 37660 41020 37716
rect 41076 37660 41086 37716
rect 57922 37660 57932 37716
rect 57988 37660 60000 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 59200 37632 60000 37660
rect 10434 37548 10444 37604
rect 10500 37548 17444 37604
rect 22978 37548 22988 37604
rect 23044 37548 26236 37604
rect 26292 37548 26572 37604
rect 26628 37548 26638 37604
rect 33506 37548 33516 37604
rect 33572 37548 35532 37604
rect 35588 37548 35598 37604
rect 15894 37436 15932 37492
rect 15988 37436 15998 37492
rect 17388 37380 17444 37548
rect 17574 37436 17612 37492
rect 17668 37436 18732 37492
rect 18788 37436 23996 37492
rect 24052 37436 24332 37492
rect 24388 37436 24398 37492
rect 27794 37436 27804 37492
rect 27860 37436 27870 37492
rect 28466 37436 28476 37492
rect 28532 37436 30716 37492
rect 30772 37436 30782 37492
rect 35634 37436 35644 37492
rect 35700 37436 36988 37492
rect 37044 37436 37054 37492
rect 37650 37436 37660 37492
rect 37716 37436 39116 37492
rect 39172 37436 39788 37492
rect 39844 37436 39854 37492
rect 44034 37436 44044 37492
rect 44100 37436 45052 37492
rect 45108 37436 45118 37492
rect 50642 37436 50652 37492
rect 50708 37436 53900 37492
rect 53956 37436 53966 37492
rect 27804 37380 27860 37436
rect 14018 37324 14028 37380
rect 14084 37324 15148 37380
rect 15204 37324 15214 37380
rect 17388 37324 23548 37380
rect 23604 37324 23614 37380
rect 25330 37324 25340 37380
rect 25396 37324 26908 37380
rect 26964 37324 26974 37380
rect 27804 37324 28588 37380
rect 28644 37324 28654 37380
rect 29250 37324 29260 37380
rect 29316 37324 29326 37380
rect 32162 37324 32172 37380
rect 32228 37324 34860 37380
rect 34916 37324 34926 37380
rect 35074 37324 35084 37380
rect 35140 37324 38108 37380
rect 38164 37324 38444 37380
rect 38500 37324 38510 37380
rect 39330 37324 39340 37380
rect 39396 37324 49756 37380
rect 49812 37324 49822 37380
rect 50372 37324 51660 37380
rect 51716 37324 51726 37380
rect 4274 37212 4284 37268
rect 4340 37212 7196 37268
rect 7252 37212 8428 37268
rect 8484 37212 9996 37268
rect 10052 37212 10062 37268
rect 10658 37212 10668 37268
rect 10724 37212 15596 37268
rect 15652 37212 15662 37268
rect 20178 37212 20188 37268
rect 20244 37212 20972 37268
rect 21028 37212 21868 37268
rect 21924 37212 21934 37268
rect 26450 37212 26460 37268
rect 26516 37212 28924 37268
rect 28980 37212 28990 37268
rect 19842 37100 19852 37156
rect 19908 37100 20524 37156
rect 20580 37100 20590 37156
rect 0 37044 800 37072
rect 29260 37044 29316 37324
rect 50372 37268 50428 37324
rect 29586 37212 29596 37268
rect 29652 37212 31948 37268
rect 32004 37212 32014 37268
rect 32274 37212 32284 37268
rect 32340 37212 33180 37268
rect 33236 37212 33246 37268
rect 44482 37212 44492 37268
rect 44548 37212 45724 37268
rect 45780 37212 45790 37268
rect 45938 37212 45948 37268
rect 46004 37212 46956 37268
rect 47012 37212 47022 37268
rect 50082 37212 50092 37268
rect 50148 37212 50428 37268
rect 50530 37212 50540 37268
rect 50596 37212 52892 37268
rect 52948 37212 52958 37268
rect 31266 37100 31276 37156
rect 31332 37100 32172 37156
rect 32228 37100 32238 37156
rect 49858 37100 49868 37156
rect 49924 37100 51436 37156
rect 51492 37100 51502 37156
rect 0 36988 2156 37044
rect 2212 36988 2222 37044
rect 27458 36988 27468 37044
rect 27524 36988 27534 37044
rect 27794 36988 27804 37044
rect 27860 36988 29316 37044
rect 30146 36988 30156 37044
rect 30212 36988 32396 37044
rect 32452 36988 32462 37044
rect 41010 36988 41020 37044
rect 41076 36988 42028 37044
rect 42084 36988 42094 37044
rect 44258 36988 44268 37044
rect 44324 36988 44940 37044
rect 44996 36988 45388 37044
rect 45444 36988 45454 37044
rect 0 36960 800 36988
rect 27468 36932 27524 36988
rect 6402 36876 6412 36932
rect 6468 36876 14588 36932
rect 14644 36876 14654 36932
rect 15362 36876 15372 36932
rect 15428 36876 16604 36932
rect 16660 36876 16670 36932
rect 21410 36876 21420 36932
rect 21476 36876 22092 36932
rect 22148 36876 24556 36932
rect 24612 36876 24622 36932
rect 27468 36876 29260 36932
rect 29316 36876 29326 36932
rect 32050 36876 32060 36932
rect 32116 36876 33068 36932
rect 33124 36876 33134 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 18274 36764 18284 36820
rect 18340 36764 18844 36820
rect 18900 36764 18910 36820
rect 29110 36764 29148 36820
rect 29204 36764 29214 36820
rect 13122 36652 13132 36708
rect 13188 36652 13916 36708
rect 13972 36652 14924 36708
rect 14980 36652 14990 36708
rect 21298 36652 21308 36708
rect 21364 36652 26236 36708
rect 26292 36652 26302 36708
rect 30370 36652 30380 36708
rect 30436 36652 32956 36708
rect 33012 36652 33022 36708
rect 34290 36652 34300 36708
rect 34356 36652 34860 36708
rect 34916 36652 35420 36708
rect 35476 36652 35486 36708
rect 36082 36652 36092 36708
rect 36148 36652 44156 36708
rect 44212 36652 44716 36708
rect 44772 36652 44782 36708
rect 46050 36652 46060 36708
rect 46116 36652 47180 36708
rect 47236 36652 47246 36708
rect 1922 36540 1932 36596
rect 1988 36540 1998 36596
rect 8978 36540 8988 36596
rect 9044 36540 11788 36596
rect 11844 36540 13468 36596
rect 13524 36540 13534 36596
rect 14476 36540 20188 36596
rect 20244 36540 20254 36596
rect 20738 36540 20748 36596
rect 20804 36540 21532 36596
rect 21588 36540 22316 36596
rect 22372 36540 22382 36596
rect 26562 36540 26572 36596
rect 26628 36540 26908 36596
rect 31490 36540 31500 36596
rect 31556 36540 41244 36596
rect 41300 36540 41804 36596
rect 41860 36540 41870 36596
rect 0 36372 800 36400
rect 1932 36372 1988 36540
rect 14476 36484 14532 36540
rect 26852 36484 26908 36540
rect 8194 36428 8204 36484
rect 8260 36428 12348 36484
rect 12404 36428 13580 36484
rect 13636 36428 13646 36484
rect 14466 36428 14476 36484
rect 14532 36428 14542 36484
rect 18946 36428 18956 36484
rect 19012 36428 19404 36484
rect 19460 36428 24052 36484
rect 26422 36428 26460 36484
rect 26516 36428 26526 36484
rect 26852 36428 27580 36484
rect 27636 36428 33964 36484
rect 34020 36428 34030 36484
rect 45266 36428 45276 36484
rect 45332 36428 46060 36484
rect 46116 36428 46126 36484
rect 23996 36372 24052 36428
rect 0 36316 1988 36372
rect 18386 36316 18396 36372
rect 18452 36316 21420 36372
rect 21476 36316 21486 36372
rect 23986 36316 23996 36372
rect 24052 36316 27356 36372
rect 27412 36316 28140 36372
rect 28196 36316 28206 36372
rect 29932 36316 30716 36372
rect 30772 36316 30782 36372
rect 30930 36316 30940 36372
rect 30996 36316 32060 36372
rect 32116 36316 32126 36372
rect 34066 36316 34076 36372
rect 34132 36316 35980 36372
rect 36036 36316 36046 36372
rect 44930 36316 44940 36372
rect 44996 36316 47292 36372
rect 47348 36316 47358 36372
rect 52994 36316 53004 36372
rect 53060 36316 54348 36372
rect 54404 36316 54414 36372
rect 0 36288 800 36316
rect 29932 36260 29988 36316
rect 7858 36204 7868 36260
rect 7924 36204 10444 36260
rect 10500 36204 10510 36260
rect 12898 36204 12908 36260
rect 12964 36204 17724 36260
rect 17780 36204 17790 36260
rect 17948 36204 23548 36260
rect 25666 36204 25676 36260
rect 25732 36204 25742 36260
rect 26674 36204 26684 36260
rect 26740 36204 29932 36260
rect 29988 36204 29998 36260
rect 39554 36204 39564 36260
rect 39620 36204 40908 36260
rect 40964 36204 42364 36260
rect 42420 36204 43036 36260
rect 43092 36204 43102 36260
rect 55346 36204 55356 36260
rect 55412 36204 56588 36260
rect 56644 36204 56654 36260
rect 17948 36148 18004 36204
rect 23492 36148 23548 36204
rect 25676 36148 25732 36204
rect 7410 36092 7420 36148
rect 7476 36092 11116 36148
rect 11172 36092 14140 36148
rect 14196 36092 14206 36148
rect 17042 36092 17052 36148
rect 17108 36092 17388 36148
rect 17444 36092 18004 36148
rect 19478 36092 19516 36148
rect 19572 36092 19582 36148
rect 23492 36092 25620 36148
rect 25676 36092 33852 36148
rect 33908 36092 35196 36148
rect 35252 36092 35262 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 25564 36036 25620 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 23314 35980 23324 36036
rect 23380 35980 23436 36036
rect 23492 35980 24668 36036
rect 24724 35980 25340 36036
rect 25396 35980 25406 36036
rect 25564 35980 26684 36036
rect 26740 35980 26750 36036
rect 27346 35980 27356 36036
rect 27412 35980 28252 36036
rect 28308 35980 28318 36036
rect 28802 35980 28812 36036
rect 28868 35980 29484 36036
rect 29540 35980 29550 36036
rect 30940 35980 34972 36036
rect 35028 35980 35038 36036
rect 14242 35868 14252 35924
rect 14308 35868 14476 35924
rect 14532 35868 14542 35924
rect 16258 35868 16268 35924
rect 16324 35868 19852 35924
rect 19908 35868 19918 35924
rect 22764 35868 23548 35924
rect 23604 35868 23614 35924
rect 24322 35868 24332 35924
rect 24388 35868 28196 35924
rect 28354 35868 28364 35924
rect 28420 35868 29372 35924
rect 29428 35868 29438 35924
rect 22764 35812 22820 35868
rect 28140 35812 28196 35868
rect 30940 35812 30996 35980
rect 34850 35868 34860 35924
rect 34916 35868 36204 35924
rect 36260 35868 36764 35924
rect 36820 35868 36830 35924
rect 43362 35868 43372 35924
rect 43428 35868 47404 35924
rect 47460 35868 47852 35924
rect 47908 35868 47918 35924
rect 13570 35756 13580 35812
rect 13636 35756 15372 35812
rect 15428 35756 15438 35812
rect 17490 35756 17500 35812
rect 17556 35756 22764 35812
rect 22820 35756 22830 35812
rect 25778 35756 25788 35812
rect 25844 35756 26908 35812
rect 28140 35756 30996 35812
rect 35858 35756 35868 35812
rect 35924 35756 37436 35812
rect 37492 35756 38108 35812
rect 38164 35756 38174 35812
rect 48066 35756 48076 35812
rect 48132 35756 49532 35812
rect 49588 35756 49598 35812
rect 0 35700 800 35728
rect 0 35644 1708 35700
rect 1764 35644 1774 35700
rect 4274 35644 4284 35700
rect 4340 35644 8988 35700
rect 9044 35644 10108 35700
rect 10164 35644 11116 35700
rect 11172 35644 11182 35700
rect 11890 35644 11900 35700
rect 11956 35644 13244 35700
rect 13300 35644 13692 35700
rect 13748 35644 13758 35700
rect 14130 35644 14140 35700
rect 14196 35644 14812 35700
rect 14868 35644 14878 35700
rect 20402 35644 20412 35700
rect 20468 35644 21308 35700
rect 21364 35644 21374 35700
rect 0 35616 800 35644
rect 11116 35588 11172 35644
rect 5506 35532 5516 35588
rect 5572 35532 6860 35588
rect 6916 35532 6926 35588
rect 11116 35532 12460 35588
rect 12516 35532 12526 35588
rect 26852 35476 26908 35756
rect 59200 35700 60000 35728
rect 27346 35644 27356 35700
rect 27412 35644 29372 35700
rect 29428 35644 29708 35700
rect 29764 35644 29774 35700
rect 34514 35644 34524 35700
rect 34580 35644 36092 35700
rect 36148 35644 36158 35700
rect 37538 35644 37548 35700
rect 37604 35644 38780 35700
rect 38836 35644 38846 35700
rect 39442 35644 39452 35700
rect 39508 35644 49084 35700
rect 49140 35644 49150 35700
rect 53218 35644 53228 35700
rect 53284 35644 53788 35700
rect 53844 35644 54236 35700
rect 54292 35644 54684 35700
rect 54740 35644 54750 35700
rect 57698 35644 57708 35700
rect 57764 35644 60000 35700
rect 59200 35616 60000 35644
rect 45714 35532 45724 35588
rect 45780 35532 46732 35588
rect 46788 35532 46798 35588
rect 26852 35420 32508 35476
rect 32564 35420 33180 35476
rect 33236 35420 33246 35476
rect 34290 35420 34300 35476
rect 34356 35420 44828 35476
rect 44884 35420 44894 35476
rect 48850 35420 48860 35476
rect 48916 35420 55804 35476
rect 55860 35420 55870 35476
rect 8530 35308 8540 35364
rect 8596 35308 9436 35364
rect 9492 35308 12012 35364
rect 12068 35308 12078 35364
rect 26338 35308 26348 35364
rect 26404 35308 34412 35364
rect 34468 35308 34478 35364
rect 35746 35308 35756 35364
rect 35812 35308 37996 35364
rect 38052 35308 38668 35364
rect 38724 35308 38734 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 14018 35196 14028 35252
rect 14084 35196 15036 35252
rect 15092 35196 16828 35252
rect 16884 35196 16894 35252
rect 19282 35196 19292 35252
rect 19348 35196 20076 35252
rect 20132 35196 29484 35252
rect 29540 35196 30044 35252
rect 30100 35196 30110 35252
rect 30258 35196 30268 35252
rect 30324 35196 31052 35252
rect 31108 35196 31118 35252
rect 37314 35196 37324 35252
rect 37380 35196 38668 35252
rect 52770 35196 52780 35252
rect 52836 35196 53340 35252
rect 53396 35196 54236 35252
rect 54292 35196 54302 35252
rect 14802 35084 14812 35140
rect 14868 35084 22260 35140
rect 22418 35084 22428 35140
rect 22484 35084 29148 35140
rect 29204 35084 29214 35140
rect 34066 35084 34076 35140
rect 34132 35084 36652 35140
rect 36708 35084 36718 35140
rect 0 35028 800 35056
rect 0 34972 1932 35028
rect 1988 34972 1998 35028
rect 8754 34972 8764 35028
rect 8820 34972 12908 35028
rect 12964 34972 13468 35028
rect 13524 34972 14476 35028
rect 14532 34972 14542 35028
rect 17826 34972 17836 35028
rect 17892 34972 19628 35028
rect 19684 34972 21980 35028
rect 22036 34972 22046 35028
rect 0 34944 800 34972
rect 8642 34860 8652 34916
rect 8708 34860 15148 34916
rect 15362 34860 15372 34916
rect 15428 34860 18620 34916
rect 18676 34860 18686 34916
rect 19394 34860 19404 34916
rect 19460 34860 21308 34916
rect 21364 34860 21374 34916
rect 8418 34748 8428 34804
rect 8484 34748 9436 34804
rect 9492 34748 11116 34804
rect 11172 34748 11182 34804
rect 15092 34692 15148 34860
rect 18620 34804 18676 34860
rect 16370 34748 16380 34804
rect 16436 34748 18396 34804
rect 18452 34748 18462 34804
rect 18620 34748 20636 34804
rect 20692 34748 20702 34804
rect 22204 34692 22260 35084
rect 38612 35028 38668 35196
rect 43026 35084 43036 35140
rect 43092 35084 47516 35140
rect 47572 35084 47582 35140
rect 49298 35084 49308 35140
rect 49364 35084 50428 35140
rect 50484 35084 50494 35140
rect 59200 35028 60000 35056
rect 22754 34972 22764 35028
rect 22820 34972 25900 35028
rect 25956 34972 26684 35028
rect 26740 34972 26750 35028
rect 32050 34972 32060 35028
rect 32116 34972 33516 35028
rect 33572 34972 33582 35028
rect 38612 34972 40572 35028
rect 40628 34972 41356 35028
rect 41412 34972 41422 35028
rect 47058 34972 47068 35028
rect 47124 34972 47628 35028
rect 47684 34972 48076 35028
rect 48132 34972 50316 35028
rect 50372 34972 50382 35028
rect 55346 34972 55356 35028
rect 55412 34972 60000 35028
rect 59200 34944 60000 34972
rect 24770 34860 24780 34916
rect 24836 34860 26348 34916
rect 26404 34860 27244 34916
rect 27300 34860 27310 34916
rect 28690 34860 28700 34916
rect 28756 34860 30940 34916
rect 30996 34860 31006 34916
rect 36306 34860 36316 34916
rect 36372 34860 37324 34916
rect 37380 34860 37390 34916
rect 46834 34860 46844 34916
rect 46900 34860 48748 34916
rect 48804 34860 48814 34916
rect 25554 34748 25564 34804
rect 25620 34748 32732 34804
rect 32788 34748 32798 34804
rect 38546 34748 38556 34804
rect 38612 34748 45164 34804
rect 45220 34748 45230 34804
rect 51986 34748 51996 34804
rect 52052 34748 52780 34804
rect 52836 34748 52846 34804
rect 54450 34748 54460 34804
rect 54516 34748 55804 34804
rect 55860 34748 55870 34804
rect 6290 34636 6300 34692
rect 6356 34636 7868 34692
rect 7924 34636 8316 34692
rect 8372 34636 8382 34692
rect 8978 34636 8988 34692
rect 9044 34636 11340 34692
rect 11396 34636 11406 34692
rect 15092 34636 21532 34692
rect 21588 34636 21598 34692
rect 22204 34636 26908 34692
rect 29474 34636 29484 34692
rect 29540 34636 30604 34692
rect 30660 34636 30670 34692
rect 43586 34636 43596 34692
rect 43652 34636 43932 34692
rect 43988 34636 43998 34692
rect 49186 34636 49196 34692
rect 49252 34636 52892 34692
rect 52948 34636 52958 34692
rect 26852 34580 26908 34636
rect 26852 34524 29932 34580
rect 29988 34524 29998 34580
rect 30146 34524 30156 34580
rect 30212 34524 34076 34580
rect 34132 34524 34142 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 5618 34412 5628 34468
rect 5684 34412 10556 34468
rect 10612 34412 14252 34468
rect 14308 34412 14700 34468
rect 14756 34412 14766 34468
rect 19030 34412 19068 34468
rect 19124 34412 19134 34468
rect 20626 34412 20636 34468
rect 20692 34412 23548 34468
rect 23604 34412 24892 34468
rect 24948 34412 24958 34468
rect 8306 34300 8316 34356
rect 8372 34300 9996 34356
rect 10052 34300 10062 34356
rect 19506 34300 19516 34356
rect 19572 34300 19852 34356
rect 19908 34300 21420 34356
rect 21476 34300 21486 34356
rect 21746 34300 21756 34356
rect 21812 34300 22988 34356
rect 23044 34300 23660 34356
rect 23716 34300 23726 34356
rect 26226 34300 26236 34356
rect 26292 34300 30380 34356
rect 30436 34300 32060 34356
rect 32116 34300 32126 34356
rect 33506 34300 33516 34356
rect 33572 34300 34188 34356
rect 34244 34300 34972 34356
rect 35028 34300 35038 34356
rect 43250 34300 43260 34356
rect 43316 34300 46508 34356
rect 46564 34300 46844 34356
rect 46900 34300 46910 34356
rect 50866 34300 50876 34356
rect 50932 34300 51436 34356
rect 51492 34300 53004 34356
rect 53060 34300 53070 34356
rect 6066 34188 6076 34244
rect 6132 34188 19628 34244
rect 19684 34188 19694 34244
rect 25666 34188 25676 34244
rect 25732 34188 30492 34244
rect 30548 34188 33628 34244
rect 33684 34188 34860 34244
rect 34916 34188 34926 34244
rect 50642 34188 50652 34244
rect 50708 34188 52444 34244
rect 52500 34188 52510 34244
rect 4834 34076 4844 34132
rect 4900 34076 5516 34132
rect 5572 34076 8316 34132
rect 8372 34076 8988 34132
rect 9044 34076 9054 34132
rect 19506 34076 19516 34132
rect 19572 34076 21532 34132
rect 21588 34076 21598 34132
rect 25554 34076 25564 34132
rect 25620 34076 26348 34132
rect 26404 34076 26414 34132
rect 32834 34076 32844 34132
rect 32900 34076 34412 34132
rect 34468 34076 34748 34132
rect 34804 34076 34814 34132
rect 50082 34076 50092 34132
rect 50148 34076 50764 34132
rect 50820 34076 50830 34132
rect 8082 33964 8092 34020
rect 8148 33964 9548 34020
rect 9604 33964 9614 34020
rect 14130 33964 14140 34020
rect 14196 33964 15260 34020
rect 15316 33964 15326 34020
rect 18386 33964 18396 34020
rect 18452 33964 24220 34020
rect 24276 33964 24286 34020
rect 3052 33852 6636 33908
rect 6692 33852 6702 33908
rect 20514 33852 20524 33908
rect 20580 33852 21308 33908
rect 21364 33852 21374 33908
rect 25666 33852 25676 33908
rect 25732 33852 26012 33908
rect 26068 33852 26078 33908
rect 36418 33852 36428 33908
rect 36484 33852 38220 33908
rect 38276 33852 38286 33908
rect 0 33684 800 33712
rect 3052 33684 3108 33852
rect 18498 33740 18508 33796
rect 18564 33740 19516 33796
rect 19572 33740 19582 33796
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 0 33628 3108 33684
rect 11106 33628 11116 33684
rect 11172 33628 13020 33684
rect 13076 33628 13412 33684
rect 0 33600 800 33628
rect 13356 33572 13412 33628
rect 39004 33628 41188 33684
rect 43922 33628 43932 33684
rect 43988 33628 45388 33684
rect 45444 33628 45454 33684
rect 39004 33572 39060 33628
rect 41132 33572 41188 33628
rect 13356 33516 14588 33572
rect 14644 33516 14654 33572
rect 18722 33516 18732 33572
rect 18788 33516 19516 33572
rect 19572 33516 19582 33572
rect 23426 33516 23436 33572
rect 23492 33516 25004 33572
rect 25060 33516 25070 33572
rect 28130 33516 28140 33572
rect 28196 33516 39060 33572
rect 39218 33516 39228 33572
rect 39284 33516 39788 33572
rect 39844 33516 40908 33572
rect 40964 33516 40974 33572
rect 41132 33516 44604 33572
rect 44660 33516 44670 33572
rect 17154 33404 17164 33460
rect 17220 33404 24332 33460
rect 24388 33404 24398 33460
rect 38210 33404 38220 33460
rect 38276 33404 38668 33460
rect 38724 33404 40460 33460
rect 40516 33404 40526 33460
rect 45948 33404 47516 33460
rect 47572 33404 47582 33460
rect 50754 33404 50764 33460
rect 50820 33404 51940 33460
rect 45948 33348 46004 33404
rect 51884 33348 51940 33404
rect 11666 33292 11676 33348
rect 11732 33292 15148 33348
rect 15250 33292 15260 33348
rect 15316 33292 16604 33348
rect 16660 33292 17500 33348
rect 17556 33292 17566 33348
rect 20402 33292 20412 33348
rect 20468 33292 20860 33348
rect 20916 33292 21980 33348
rect 22036 33292 25676 33348
rect 25732 33292 25742 33348
rect 34290 33292 34300 33348
rect 34356 33292 42476 33348
rect 42532 33292 42542 33348
rect 45266 33292 45276 33348
rect 45332 33292 45948 33348
rect 46004 33292 46014 33348
rect 47170 33292 47180 33348
rect 47236 33292 48636 33348
rect 48692 33292 49532 33348
rect 49588 33292 49598 33348
rect 50194 33292 50204 33348
rect 50260 33292 50876 33348
rect 50932 33292 50942 33348
rect 51874 33292 51884 33348
rect 51940 33292 53004 33348
rect 53060 33292 53070 33348
rect 54338 33292 54348 33348
rect 54404 33292 55580 33348
rect 55636 33292 55646 33348
rect 15092 33236 15148 33292
rect 2034 33180 2044 33236
rect 2100 33180 7532 33236
rect 7588 33180 7598 33236
rect 13682 33180 13692 33236
rect 13748 33180 14420 33236
rect 15092 33180 22092 33236
rect 22148 33180 22158 33236
rect 24434 33180 24444 33236
rect 24500 33180 25564 33236
rect 25620 33180 27020 33236
rect 27076 33180 27086 33236
rect 43138 33180 43148 33236
rect 43204 33180 43596 33236
rect 43652 33180 43662 33236
rect 45602 33180 45612 33236
rect 45668 33180 46284 33236
rect 46340 33180 47068 33236
rect 47124 33180 48188 33236
rect 48244 33180 48254 33236
rect 48514 33180 48524 33236
rect 48580 33180 51324 33236
rect 51380 33180 51390 33236
rect 14364 33124 14420 33180
rect 12002 33068 12012 33124
rect 12068 33068 12572 33124
rect 12628 33068 13580 33124
rect 13636 33068 14028 33124
rect 14084 33068 14094 33124
rect 14364 33068 18956 33124
rect 19012 33068 19022 33124
rect 19628 33068 23996 33124
rect 24052 33068 24780 33124
rect 24836 33068 25452 33124
rect 25508 33068 25900 33124
rect 25956 33068 25966 33124
rect 50082 33068 50092 33124
rect 50148 33068 51436 33124
rect 51492 33068 51502 33124
rect 0 33012 800 33040
rect 19628 33012 19684 33068
rect 59200 33012 60000 33040
rect 0 32956 1708 33012
rect 1764 32956 2492 33012
rect 2548 32956 2558 33012
rect 19058 32956 19068 33012
rect 19124 32956 19684 33012
rect 37538 32956 37548 33012
rect 37604 32956 43148 33012
rect 43204 32956 43708 33012
rect 43764 32956 43774 33012
rect 57922 32956 57932 33012
rect 57988 32956 60000 33012
rect 0 32928 800 32956
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 59200 32928 60000 32956
rect 19142 32844 19180 32900
rect 19236 32844 19246 32900
rect 10882 32732 10892 32788
rect 10948 32732 28588 32788
rect 28644 32732 29484 32788
rect 29540 32732 29550 32788
rect 29810 32732 29820 32788
rect 29876 32732 31724 32788
rect 31780 32732 31790 32788
rect 36194 32732 36204 32788
rect 36260 32732 37212 32788
rect 37268 32732 38108 32788
rect 38164 32732 38174 32788
rect 47506 32732 47516 32788
rect 47572 32732 48076 32788
rect 48132 32732 49196 32788
rect 49252 32732 49644 32788
rect 49700 32732 49710 32788
rect 18498 32620 18508 32676
rect 18564 32620 19852 32676
rect 19908 32620 23436 32676
rect 23492 32620 25228 32676
rect 25284 32620 26908 32676
rect 26964 32620 26974 32676
rect 36642 32620 36652 32676
rect 36708 32620 37324 32676
rect 37380 32620 37772 32676
rect 37828 32620 37838 32676
rect 43922 32620 43932 32676
rect 43988 32620 46956 32676
rect 47012 32620 47628 32676
rect 47684 32620 47694 32676
rect 30146 32508 30156 32564
rect 30212 32508 30828 32564
rect 30884 32508 37212 32564
rect 37268 32508 37548 32564
rect 37604 32508 37614 32564
rect 49522 32508 49532 32564
rect 49588 32508 49868 32564
rect 49924 32508 49934 32564
rect 29250 32396 29260 32452
rect 29316 32396 30604 32452
rect 30660 32396 30670 32452
rect 23090 32284 23100 32340
rect 23156 32284 23548 32340
rect 23604 32284 24220 32340
rect 24276 32284 24286 32340
rect 41010 32172 41020 32228
rect 41076 32172 42700 32228
rect 42756 32172 42766 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 30818 31948 30828 32004
rect 30884 31948 32732 32004
rect 32788 31948 32798 32004
rect 48178 31948 48188 32004
rect 48244 31948 48860 32004
rect 48916 31948 48926 32004
rect 21186 31836 21196 31892
rect 21252 31836 31388 31892
rect 31444 31836 31454 31892
rect 32172 31836 42868 31892
rect 43026 31836 43036 31892
rect 43092 31836 43708 31892
rect 43764 31836 44156 31892
rect 44212 31836 44222 31892
rect 32172 31780 32228 31836
rect 42812 31780 42868 31836
rect 10098 31724 10108 31780
rect 10164 31724 21980 31780
rect 22036 31724 22046 31780
rect 25218 31724 25228 31780
rect 25284 31724 26124 31780
rect 26180 31724 26190 31780
rect 28466 31724 28476 31780
rect 28532 31724 32228 31780
rect 34178 31724 34188 31780
rect 34244 31724 38668 31780
rect 38724 31724 38734 31780
rect 42812 31724 44044 31780
rect 44100 31724 44110 31780
rect 0 31668 800 31696
rect 0 31612 2380 31668
rect 2436 31612 2446 31668
rect 0 31584 800 31612
rect 2034 31500 2044 31556
rect 2100 31500 17500 31556
rect 17556 31500 18172 31556
rect 18228 31500 18238 31556
rect 19954 31500 19964 31556
rect 20020 31500 25788 31556
rect 25844 31500 25854 31556
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 26124 31332 26180 31724
rect 32946 31612 32956 31668
rect 33012 31612 33740 31668
rect 33796 31612 33806 31668
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 20188 31276 26068 31332
rect 26124 31276 28140 31332
rect 28196 31276 30044 31332
rect 30100 31276 31836 31332
rect 31892 31276 33180 31332
rect 33236 31276 33628 31332
rect 33684 31276 33694 31332
rect 20188 31220 20244 31276
rect 26012 31220 26068 31276
rect 17826 31164 17836 31220
rect 17892 31164 18956 31220
rect 19012 31164 19022 31220
rect 19170 31164 19180 31220
rect 19236 31164 20244 31220
rect 25778 31164 25788 31220
rect 25844 31164 25854 31220
rect 26012 31164 36540 31220
rect 36596 31164 36606 31220
rect 38322 31164 38332 31220
rect 38388 31164 38780 31220
rect 38836 31164 38846 31220
rect 38994 31164 39004 31220
rect 39060 31164 41692 31220
rect 41748 31164 41758 31220
rect 41906 31164 41916 31220
rect 41972 31164 45388 31220
rect 45444 31164 45454 31220
rect 25788 31108 25844 31164
rect 16706 31052 16716 31108
rect 16772 31052 21868 31108
rect 21924 31052 21934 31108
rect 25788 31052 31948 31108
rect 32004 31052 32956 31108
rect 33012 31052 33628 31108
rect 33684 31052 33694 31108
rect 33954 31052 33964 31108
rect 34020 31052 57820 31108
rect 57876 31052 57886 31108
rect 0 30996 800 31024
rect 21868 30996 21924 31052
rect 0 30940 1820 30996
rect 1876 30940 1886 30996
rect 6626 30940 6636 30996
rect 6692 30940 18956 30996
rect 19012 30940 19404 30996
rect 19460 30940 19470 30996
rect 21868 30940 26908 30996
rect 26964 30940 26974 30996
rect 39778 30940 39788 30996
rect 39844 30940 41356 30996
rect 41412 30940 41422 30996
rect 0 30912 800 30940
rect 21746 30828 21756 30884
rect 21812 30828 24444 30884
rect 24500 30828 24510 30884
rect 25554 30828 25564 30884
rect 25620 30828 25900 30884
rect 25956 30828 26236 30884
rect 26292 30828 26572 30884
rect 26628 30828 26638 30884
rect 40338 30828 40348 30884
rect 40404 30828 41020 30884
rect 41076 30828 41086 30884
rect 4274 30716 4284 30772
rect 4340 30716 21308 30772
rect 21364 30716 23996 30772
rect 24052 30716 24062 30772
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 17042 30492 17052 30548
rect 17108 30492 28700 30548
rect 28756 30492 28766 30548
rect 13906 30380 13916 30436
rect 13972 30380 15484 30436
rect 15540 30380 15550 30436
rect 19170 30380 19180 30436
rect 19236 30380 20076 30436
rect 20132 30380 20142 30436
rect 38882 30380 38892 30436
rect 38948 30380 39676 30436
rect 39732 30380 39742 30436
rect 0 30324 800 30352
rect 59200 30324 60000 30352
rect 0 30268 1932 30324
rect 1988 30268 1998 30324
rect 11666 30268 11676 30324
rect 11732 30268 27804 30324
rect 27860 30268 27870 30324
rect 58146 30268 58156 30324
rect 58212 30268 60000 30324
rect 0 30240 800 30268
rect 59200 30240 60000 30268
rect 8754 30156 8764 30212
rect 8820 30156 11228 30212
rect 11284 30156 11788 30212
rect 11844 30156 11854 30212
rect 13682 30156 13692 30212
rect 13748 30156 19404 30212
rect 19460 30156 19470 30212
rect 20066 30156 20076 30212
rect 20132 30156 22316 30212
rect 22372 30156 22382 30212
rect 23762 30156 23772 30212
rect 23828 30156 24668 30212
rect 24724 30156 24734 30212
rect 31826 30156 31836 30212
rect 31892 30156 32060 30212
rect 32116 30156 32620 30212
rect 32676 30156 33964 30212
rect 34020 30156 34030 30212
rect 5954 30044 5964 30100
rect 6020 30044 6030 30100
rect 7858 30044 7868 30100
rect 7924 30044 8540 30100
rect 8596 30044 8606 30100
rect 9874 30044 9884 30100
rect 9940 30044 10780 30100
rect 10836 30044 10846 30100
rect 15092 30044 16940 30100
rect 16996 30044 17006 30100
rect 19282 30044 19292 30100
rect 19348 30044 21308 30100
rect 21364 30044 21374 30100
rect 32722 30044 32732 30100
rect 32788 30044 33292 30100
rect 33348 30044 33358 30100
rect 44258 30044 44268 30100
rect 44324 30044 45612 30100
rect 45668 30044 45678 30100
rect 5964 29988 6020 30044
rect 15092 29988 15148 30044
rect 5964 29932 15148 29988
rect 21746 29932 21756 29988
rect 21812 29932 22540 29988
rect 22596 29932 22606 29988
rect 24322 29932 24332 29988
rect 24388 29932 25676 29988
rect 25732 29932 25742 29988
rect 27906 29932 27916 29988
rect 27972 29932 30828 29988
rect 30884 29932 30894 29988
rect 38546 29932 38556 29988
rect 38612 29932 39228 29988
rect 39284 29932 39294 29988
rect 7186 29820 7196 29876
rect 7252 29820 9100 29876
rect 9156 29820 9166 29876
rect 20626 29820 20636 29876
rect 20692 29820 30268 29876
rect 30324 29820 30334 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 0 29652 800 29680
rect 0 29596 2492 29652
rect 2548 29596 2558 29652
rect 17714 29596 17724 29652
rect 17780 29596 19964 29652
rect 20020 29596 20636 29652
rect 20692 29596 21196 29652
rect 21252 29596 21262 29652
rect 21970 29596 21980 29652
rect 22036 29596 23996 29652
rect 24052 29596 25116 29652
rect 25172 29596 25182 29652
rect 31602 29596 31612 29652
rect 31668 29596 32172 29652
rect 32228 29596 33404 29652
rect 33460 29596 33470 29652
rect 36306 29596 36316 29652
rect 36372 29596 37324 29652
rect 37380 29596 37390 29652
rect 38434 29596 38444 29652
rect 38500 29596 39452 29652
rect 39508 29596 39518 29652
rect 0 29568 800 29596
rect 11004 29484 17500 29540
rect 17556 29484 17948 29540
rect 18004 29484 18014 29540
rect 19842 29484 19852 29540
rect 19908 29484 22204 29540
rect 22260 29484 22270 29540
rect 24658 29484 24668 29540
rect 24724 29484 25452 29540
rect 25508 29484 26236 29540
rect 26292 29484 27580 29540
rect 27636 29484 27646 29540
rect 11004 29428 11060 29484
rect 10994 29372 11004 29428
rect 11060 29372 11070 29428
rect 14354 29372 14364 29428
rect 14420 29372 15372 29428
rect 15428 29372 15438 29428
rect 15586 29372 15596 29428
rect 15652 29372 15662 29428
rect 17602 29372 17612 29428
rect 17668 29372 17836 29428
rect 17892 29372 17902 29428
rect 18050 29372 18060 29428
rect 18116 29372 19796 29428
rect 28578 29372 28588 29428
rect 28644 29372 29148 29428
rect 29204 29372 29214 29428
rect 33058 29372 33068 29428
rect 33124 29372 33740 29428
rect 33796 29372 33806 29428
rect 43250 29372 43260 29428
rect 43316 29372 43932 29428
rect 43988 29372 43998 29428
rect 15596 29316 15652 29372
rect 19740 29316 19796 29372
rect 9762 29260 9772 29316
rect 9828 29260 10444 29316
rect 10500 29260 10510 29316
rect 15092 29260 15652 29316
rect 16678 29260 16716 29316
rect 16772 29260 16782 29316
rect 18946 29260 18956 29316
rect 19012 29260 19022 29316
rect 19730 29260 19740 29316
rect 19796 29260 20748 29316
rect 20804 29260 20814 29316
rect 21298 29260 21308 29316
rect 21364 29260 21644 29316
rect 21700 29260 22876 29316
rect 22932 29260 22942 29316
rect 26852 29260 39116 29316
rect 39172 29260 39564 29316
rect 39620 29260 40236 29316
rect 40292 29260 40302 29316
rect 15092 29204 15148 29260
rect 1922 29148 1932 29204
rect 1988 29148 1998 29204
rect 10994 29148 11004 29204
rect 11060 29148 12460 29204
rect 12516 29148 15148 29204
rect 18498 29148 18508 29204
rect 18564 29148 18732 29204
rect 18788 29148 18798 29204
rect 0 28980 800 29008
rect 1932 28980 1988 29148
rect 18956 29092 19012 29260
rect 5058 29036 5068 29092
rect 5124 29036 19012 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 0 28924 1988 28980
rect 10994 28924 11004 28980
rect 11060 28924 15148 28980
rect 18610 28924 18620 28980
rect 18676 28924 19348 28980
rect 0 28896 800 28924
rect 15092 28868 15148 28924
rect 19292 28868 19348 28924
rect 26852 28868 26908 29260
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 4274 28812 4284 28868
rect 4340 28812 12012 28868
rect 12068 28812 13468 28868
rect 13524 28812 13534 28868
rect 15092 28812 18452 28868
rect 19282 28812 19292 28868
rect 19348 28812 26908 28868
rect 33282 28812 33292 28868
rect 33348 28812 37604 28868
rect 13468 28756 13524 28812
rect 18396 28756 18452 28812
rect 5954 28700 5964 28756
rect 6020 28700 7756 28756
rect 7812 28700 10556 28756
rect 10612 28700 10622 28756
rect 13468 28700 16044 28756
rect 16100 28700 16380 28756
rect 16436 28700 16446 28756
rect 18396 28700 21700 28756
rect 21970 28700 21980 28756
rect 22036 28700 31948 28756
rect 32004 28700 32014 28756
rect 33170 28700 33180 28756
rect 33236 28700 33964 28756
rect 34020 28700 37324 28756
rect 37380 28700 37390 28756
rect 21644 28644 21700 28700
rect 31948 28644 32004 28700
rect 37548 28644 37604 28812
rect 4274 28588 4284 28644
rect 4340 28588 6972 28644
rect 7028 28588 7644 28644
rect 7700 28588 7710 28644
rect 9202 28588 9212 28644
rect 9268 28588 10108 28644
rect 10164 28588 10174 28644
rect 13906 28588 13916 28644
rect 13972 28588 14700 28644
rect 14756 28588 15484 28644
rect 15540 28588 15550 28644
rect 17602 28588 17612 28644
rect 17668 28588 19740 28644
rect 19796 28588 20524 28644
rect 20580 28588 20590 28644
rect 21634 28588 21644 28644
rect 21700 28588 21710 28644
rect 22754 28588 22764 28644
rect 22820 28588 26124 28644
rect 26180 28588 26190 28644
rect 29474 28588 29484 28644
rect 29540 28588 31052 28644
rect 31108 28588 31118 28644
rect 31948 28588 34972 28644
rect 35028 28588 35252 28644
rect 35634 28588 35644 28644
rect 35700 28588 37212 28644
rect 37268 28588 37278 28644
rect 37538 28588 37548 28644
rect 37604 28588 38220 28644
rect 38276 28588 38286 28644
rect 35196 28532 35252 28588
rect 4162 28476 4172 28532
rect 4228 28476 6636 28532
rect 6692 28476 8428 28532
rect 8484 28476 8494 28532
rect 15586 28476 15596 28532
rect 15652 28476 16716 28532
rect 16772 28476 18956 28532
rect 19012 28476 24668 28532
rect 24724 28476 24734 28532
rect 35196 28476 35532 28532
rect 35588 28476 35598 28532
rect 37090 28476 37100 28532
rect 37156 28476 38332 28532
rect 38388 28476 38398 28532
rect 9090 28364 9100 28420
rect 9156 28364 20300 28420
rect 20356 28364 21532 28420
rect 21588 28364 21598 28420
rect 22306 28364 22316 28420
rect 22372 28364 23100 28420
rect 23156 28364 23166 28420
rect 31266 28364 31276 28420
rect 31332 28364 32956 28420
rect 33012 28364 38780 28420
rect 38836 28364 39788 28420
rect 39844 28364 39854 28420
rect 0 28308 800 28336
rect 59200 28308 60000 28336
rect 0 28252 1932 28308
rect 1988 28252 1998 28308
rect 20626 28252 20636 28308
rect 20692 28252 32396 28308
rect 32452 28252 32462 28308
rect 58146 28252 58156 28308
rect 58212 28252 60000 28308
rect 0 28224 800 28252
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 59200 28224 60000 28252
rect 16258 28028 16268 28084
rect 16324 28028 22764 28084
rect 22820 28028 22830 28084
rect 24658 28028 24668 28084
rect 24724 28028 25676 28084
rect 25732 28028 26124 28084
rect 26180 28028 26908 28084
rect 26964 28028 26974 28084
rect 27682 28028 27692 28084
rect 27748 28028 28588 28084
rect 28644 28028 29036 28084
rect 29092 28028 29820 28084
rect 29876 28028 29886 28084
rect 30930 28028 30940 28084
rect 30996 28028 33964 28084
rect 34020 28028 34030 28084
rect 42578 28028 42588 28084
rect 42644 28028 43932 28084
rect 43988 28028 45164 28084
rect 45220 28028 45612 28084
rect 45668 28028 45678 28084
rect 8418 27916 8428 27972
rect 8484 27916 9548 27972
rect 9604 27916 9614 27972
rect 9874 27916 9884 27972
rect 9940 27916 10892 27972
rect 10948 27916 11228 27972
rect 11284 27916 12348 27972
rect 12404 27916 12414 27972
rect 15138 27916 15148 27972
rect 15204 27916 16268 27972
rect 16324 27916 16334 27972
rect 16930 27916 16940 27972
rect 16996 27916 17612 27972
rect 17668 27916 22316 27972
rect 22372 27916 22382 27972
rect 36866 27916 36876 27972
rect 36932 27916 41356 27972
rect 41412 27916 41422 27972
rect 9762 27804 9772 27860
rect 9828 27804 10780 27860
rect 10836 27804 10846 27860
rect 14018 27804 14028 27860
rect 14084 27804 17388 27860
rect 17444 27804 17454 27860
rect 22530 27804 22540 27860
rect 22596 27804 27468 27860
rect 27524 27804 27534 27860
rect 39778 27804 39788 27860
rect 39844 27804 40796 27860
rect 40852 27804 40862 27860
rect 14354 27692 14364 27748
rect 14420 27692 17780 27748
rect 17938 27692 17948 27748
rect 18004 27692 19404 27748
rect 19460 27692 19470 27748
rect 27794 27692 27804 27748
rect 27860 27692 28252 27748
rect 28308 27692 28318 27748
rect 0 27636 800 27664
rect 17724 27636 17780 27692
rect 0 27580 1932 27636
rect 1988 27580 1998 27636
rect 7298 27580 7308 27636
rect 7364 27580 8092 27636
rect 8148 27580 8158 27636
rect 11666 27580 11676 27636
rect 11732 27580 15148 27636
rect 17724 27580 28924 27636
rect 28980 27580 28990 27636
rect 35522 27580 35532 27636
rect 35588 27580 37436 27636
rect 37492 27580 37502 27636
rect 38612 27580 44492 27636
rect 44548 27580 44558 27636
rect 0 27552 800 27580
rect 15092 27524 15148 27580
rect 38612 27524 38668 27580
rect 11218 27468 11228 27524
rect 11284 27468 14028 27524
rect 14084 27468 14094 27524
rect 15092 27468 23548 27524
rect 23604 27468 23614 27524
rect 25442 27468 25452 27524
rect 25508 27468 28476 27524
rect 28532 27468 28542 27524
rect 35746 27468 35756 27524
rect 35812 27468 38668 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 10434 27356 10444 27412
rect 10500 27356 11004 27412
rect 11060 27356 15764 27412
rect 16818 27356 16828 27412
rect 16884 27356 19852 27412
rect 19908 27356 21532 27412
rect 21588 27356 21598 27412
rect 8530 27244 8540 27300
rect 8596 27244 11116 27300
rect 11172 27244 13244 27300
rect 13300 27244 13804 27300
rect 13860 27244 13870 27300
rect 9538 27132 9548 27188
rect 9604 27132 12236 27188
rect 12292 27132 12302 27188
rect 14242 27132 14252 27188
rect 14308 27132 14700 27188
rect 14756 27132 14766 27188
rect 15708 27076 15764 27356
rect 16258 27244 16268 27300
rect 16324 27244 18564 27300
rect 18508 27188 18564 27244
rect 16594 27132 16604 27188
rect 16660 27132 17612 27188
rect 17668 27132 17678 27188
rect 18498 27132 18508 27188
rect 18564 27132 18574 27188
rect 22754 27132 22764 27188
rect 22820 27132 26236 27188
rect 26292 27132 26302 27188
rect 31714 27132 31724 27188
rect 31780 27132 32284 27188
rect 32340 27132 35756 27188
rect 35812 27132 35822 27188
rect 36418 27132 36428 27188
rect 36484 27132 37100 27188
rect 37156 27132 37166 27188
rect 41458 27132 41468 27188
rect 41524 27132 42588 27188
rect 42644 27132 42654 27188
rect 6066 27020 6076 27076
rect 6132 27020 7308 27076
rect 7364 27020 7374 27076
rect 7522 27020 7532 27076
rect 7588 27020 10444 27076
rect 10500 27020 10510 27076
rect 10882 27020 10892 27076
rect 10948 27020 11564 27076
rect 11620 27020 11630 27076
rect 12898 27020 12908 27076
rect 12964 27020 15148 27076
rect 15698 27020 15708 27076
rect 15764 27020 18060 27076
rect 18116 27020 18126 27076
rect 26450 27020 26460 27076
rect 26516 27020 27132 27076
rect 27188 27020 27804 27076
rect 27860 27020 29148 27076
rect 29204 27020 29214 27076
rect 34962 27020 34972 27076
rect 35028 27020 36988 27076
rect 37044 27020 37054 27076
rect 39218 27020 39228 27076
rect 39284 27020 42364 27076
rect 42420 27020 43484 27076
rect 43540 27020 43550 27076
rect 0 26964 800 26992
rect 15092 26964 15148 27020
rect 0 26908 1708 26964
rect 1764 26908 1774 26964
rect 4834 26908 4844 26964
rect 4900 26908 8988 26964
rect 9044 26908 9054 26964
rect 12114 26908 12124 26964
rect 12180 26908 13356 26964
rect 13412 26908 13692 26964
rect 13748 26908 13758 26964
rect 15092 26908 16268 26964
rect 16324 26908 16334 26964
rect 16828 26908 21308 26964
rect 21364 26908 21374 26964
rect 23314 26908 23324 26964
rect 23380 26908 25788 26964
rect 25844 26908 25854 26964
rect 28802 26908 28812 26964
rect 28868 26908 29260 26964
rect 29316 26908 29326 26964
rect 0 26880 800 26908
rect 16828 26740 16884 26908
rect 17826 26796 17836 26852
rect 17892 26796 20748 26852
rect 20804 26796 20814 26852
rect 24322 26796 24332 26852
rect 24388 26796 27244 26852
rect 27300 26796 28588 26852
rect 28644 26796 28654 26852
rect 12450 26684 12460 26740
rect 12516 26684 13916 26740
rect 13972 26684 13982 26740
rect 14242 26684 14252 26740
rect 14308 26684 16884 26740
rect 19366 26684 19404 26740
rect 19460 26684 19470 26740
rect 19618 26684 19628 26740
rect 19684 26684 19694 26740
rect 19628 26628 19684 26684
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 15362 26572 15372 26628
rect 15428 26572 18732 26628
rect 18788 26572 19684 26628
rect 13458 26460 13468 26516
rect 13524 26460 13916 26516
rect 13972 26460 18676 26516
rect 19394 26460 19404 26516
rect 19460 26460 22988 26516
rect 23044 26460 23054 26516
rect 18620 26292 18676 26460
rect 19842 26348 19852 26404
rect 19908 26348 20524 26404
rect 20580 26348 20590 26404
rect 20850 26348 20860 26404
rect 20916 26348 24780 26404
rect 24836 26348 24846 26404
rect 59200 26292 60000 26320
rect 9426 26236 9436 26292
rect 9492 26236 10108 26292
rect 10164 26236 10668 26292
rect 10724 26236 10734 26292
rect 13570 26236 13580 26292
rect 13636 26236 15260 26292
rect 15316 26236 15326 26292
rect 16146 26236 16156 26292
rect 16212 26236 16716 26292
rect 16772 26236 16782 26292
rect 17378 26236 17388 26292
rect 17444 26236 18172 26292
rect 18228 26236 18238 26292
rect 18610 26236 18620 26292
rect 18676 26236 18686 26292
rect 18834 26236 18844 26292
rect 18900 26236 19740 26292
rect 19796 26236 19806 26292
rect 20178 26236 20188 26292
rect 20244 26236 21756 26292
rect 21812 26236 21822 26292
rect 29362 26236 29372 26292
rect 29428 26236 30380 26292
rect 30436 26236 30446 26292
rect 39218 26236 39228 26292
rect 39284 26236 42252 26292
rect 42308 26236 42318 26292
rect 58258 26236 58268 26292
rect 58324 26236 60000 26292
rect 59200 26208 60000 26236
rect 6850 26124 6860 26180
rect 6916 26124 13020 26180
rect 13076 26124 13468 26180
rect 13524 26124 14364 26180
rect 14420 26124 14430 26180
rect 16370 26124 16380 26180
rect 16436 26124 16828 26180
rect 16884 26124 18060 26180
rect 18116 26124 18126 26180
rect 18274 26124 18284 26180
rect 18340 26124 19068 26180
rect 19124 26124 19134 26180
rect 20402 26124 20412 26180
rect 20468 26124 24332 26180
rect 24388 26124 24398 26180
rect 20412 26068 20468 26124
rect 7410 26012 7420 26068
rect 7476 26012 14252 26068
rect 14308 26012 14318 26068
rect 14476 26012 15596 26068
rect 15652 26012 15662 26068
rect 17378 26012 17388 26068
rect 17444 26012 20468 26068
rect 23986 26012 23996 26068
rect 24052 26012 25788 26068
rect 25844 26012 25854 26068
rect 27346 26012 27356 26068
rect 27412 26012 28476 26068
rect 28532 26012 30716 26068
rect 30772 26012 31052 26068
rect 31108 26012 31118 26068
rect 43474 26012 43484 26068
rect 43540 26012 45948 26068
rect 46004 26012 46014 26068
rect 14476 25956 14532 26012
rect 12114 25900 12124 25956
rect 12180 25900 13692 25956
rect 13748 25900 14532 25956
rect 14802 25900 14812 25956
rect 14868 25900 15372 25956
rect 15428 25900 15438 25956
rect 16044 25900 17500 25956
rect 17556 25900 17566 25956
rect 22194 25900 22204 25956
rect 22260 25900 23436 25956
rect 23492 25900 26012 25956
rect 26068 25900 26078 25956
rect 27906 25900 27916 25956
rect 27972 25900 28140 25956
rect 28196 25900 30268 25956
rect 30324 25900 31276 25956
rect 31332 25900 31342 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 16044 25844 16100 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 6402 25788 6412 25844
rect 6468 25788 14140 25844
rect 14196 25788 14206 25844
rect 14354 25788 14364 25844
rect 14420 25788 16100 25844
rect 16258 25788 16268 25844
rect 16324 25788 25228 25844
rect 25284 25788 25294 25844
rect 29138 25788 29148 25844
rect 29204 25788 29708 25844
rect 29764 25788 29774 25844
rect 9314 25676 9324 25732
rect 9380 25676 10556 25732
rect 10612 25676 10622 25732
rect 11890 25676 11900 25732
rect 11956 25676 14476 25732
rect 14532 25676 14542 25732
rect 15092 25676 19852 25732
rect 19908 25676 19918 25732
rect 20850 25676 20860 25732
rect 20916 25676 32060 25732
rect 32116 25676 32126 25732
rect 0 25620 800 25648
rect 0 25564 2156 25620
rect 2212 25564 2222 25620
rect 11666 25564 11676 25620
rect 11732 25564 13804 25620
rect 13860 25564 13870 25620
rect 14354 25564 14364 25620
rect 14420 25564 14812 25620
rect 14868 25564 14878 25620
rect 0 25536 800 25564
rect 15092 25508 15148 25676
rect 59200 25620 60000 25648
rect 17826 25564 17836 25620
rect 17892 25564 18172 25620
rect 18228 25564 18238 25620
rect 19506 25564 19516 25620
rect 19572 25564 29148 25620
rect 29204 25564 29932 25620
rect 29988 25564 29998 25620
rect 32162 25564 32172 25620
rect 32228 25564 35196 25620
rect 35252 25564 36092 25620
rect 36148 25564 36158 25620
rect 58146 25564 58156 25620
rect 58212 25564 60000 25620
rect 59200 25536 60000 25564
rect 5954 25452 5964 25508
rect 6020 25452 8092 25508
rect 8148 25452 8158 25508
rect 8642 25452 8652 25508
rect 8708 25452 9324 25508
rect 9380 25452 9884 25508
rect 9940 25452 9950 25508
rect 10994 25452 11004 25508
rect 11060 25452 11452 25508
rect 11508 25452 12236 25508
rect 12292 25452 12302 25508
rect 12674 25452 12684 25508
rect 12740 25452 13916 25508
rect 13972 25452 13982 25508
rect 14242 25452 14252 25508
rect 14308 25452 15148 25508
rect 15362 25452 15372 25508
rect 15428 25452 15932 25508
rect 15988 25452 15998 25508
rect 17490 25452 17500 25508
rect 17556 25452 20188 25508
rect 20244 25452 20254 25508
rect 22306 25452 22316 25508
rect 22372 25452 23212 25508
rect 23268 25452 23884 25508
rect 23940 25452 23950 25508
rect 25106 25452 25116 25508
rect 25172 25452 28252 25508
rect 28308 25452 28318 25508
rect 28578 25452 28588 25508
rect 28644 25452 30044 25508
rect 30100 25452 30110 25508
rect 43362 25452 43372 25508
rect 43428 25452 43932 25508
rect 43988 25452 43998 25508
rect 47058 25452 47068 25508
rect 47124 25452 55580 25508
rect 55636 25452 55646 25508
rect 5618 25340 5628 25396
rect 5684 25340 6860 25396
rect 6916 25340 6926 25396
rect 11330 25340 11340 25396
rect 11396 25340 11788 25396
rect 11844 25340 11854 25396
rect 12012 25340 12460 25396
rect 12516 25340 12526 25396
rect 13010 25340 13020 25396
rect 13076 25340 17724 25396
rect 17780 25340 17790 25396
rect 21522 25340 21532 25396
rect 21588 25340 26124 25396
rect 26180 25340 26190 25396
rect 27570 25340 27580 25396
rect 27636 25340 27916 25396
rect 27972 25340 27982 25396
rect 28354 25340 28364 25396
rect 28420 25340 29260 25396
rect 29316 25340 29326 25396
rect 12012 25284 12068 25340
rect 9874 25228 9884 25284
rect 9940 25228 12012 25284
rect 12068 25228 12078 25284
rect 16482 25228 16492 25284
rect 16548 25228 17836 25284
rect 17892 25228 17902 25284
rect 21420 25228 21756 25284
rect 21812 25228 22540 25284
rect 22596 25228 22606 25284
rect 24658 25228 24668 25284
rect 24724 25228 25340 25284
rect 25396 25228 27692 25284
rect 27748 25228 27758 25284
rect 31798 25228 31836 25284
rect 31892 25228 31902 25284
rect 36194 25228 36204 25284
rect 36260 25228 36988 25284
rect 37044 25228 37884 25284
rect 37940 25228 37950 25284
rect 42690 25228 42700 25284
rect 42756 25228 43484 25284
rect 43540 25228 43550 25284
rect 8978 25116 8988 25172
rect 9044 25116 14812 25172
rect 14868 25116 14878 25172
rect 15026 25116 15036 25172
rect 15092 25116 15820 25172
rect 15876 25116 15886 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 13570 25004 13580 25060
rect 13636 25004 14700 25060
rect 14756 25004 15708 25060
rect 15764 25004 15774 25060
rect 11890 24892 11900 24948
rect 11956 24892 12908 24948
rect 12964 24892 13468 24948
rect 13524 24892 14140 24948
rect 14196 24892 14206 24948
rect 14588 24892 16268 24948
rect 16324 24892 16334 24948
rect 14588 24836 14644 24892
rect 21420 24836 21476 25228
rect 28242 25116 28252 25172
rect 28308 25116 28476 25172
rect 28532 25116 29596 25172
rect 29652 25116 30604 25172
rect 30660 25116 30670 25172
rect 42802 25116 42812 25172
rect 42868 25116 44828 25172
rect 44884 25116 44894 25172
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 59200 24948 60000 24976
rect 22306 24892 22316 24948
rect 22372 24892 23212 24948
rect 23268 24892 23278 24948
rect 25218 24892 25228 24948
rect 25284 24892 30604 24948
rect 30660 24892 30670 24948
rect 37314 24892 37324 24948
rect 37380 24892 38892 24948
rect 38948 24892 38958 24948
rect 57922 24892 57932 24948
rect 57988 24892 60000 24948
rect 59200 24864 60000 24892
rect 8978 24780 8988 24836
rect 9044 24780 11452 24836
rect 11508 24780 11518 24836
rect 13010 24780 13020 24836
rect 13076 24780 14644 24836
rect 14924 24780 16716 24836
rect 16772 24780 16782 24836
rect 19394 24780 19404 24836
rect 19460 24780 20972 24836
rect 21028 24780 21038 24836
rect 21410 24780 21420 24836
rect 21476 24780 21486 24836
rect 28662 24780 28700 24836
rect 28756 24780 28766 24836
rect 30146 24780 30156 24836
rect 30212 24780 31164 24836
rect 31220 24780 31230 24836
rect 41346 24780 41356 24836
rect 41412 24780 43260 24836
rect 43316 24780 43326 24836
rect 7858 24668 7868 24724
rect 7924 24668 8540 24724
rect 8596 24668 9548 24724
rect 9604 24668 9614 24724
rect 14924 24612 14980 24780
rect 17714 24668 17724 24724
rect 17780 24668 20188 24724
rect 20244 24668 20254 24724
rect 20748 24668 25340 24724
rect 25396 24668 25564 24724
rect 25620 24668 25630 24724
rect 31826 24668 31836 24724
rect 31892 24668 33180 24724
rect 33236 24668 33852 24724
rect 33908 24668 33918 24724
rect 20748 24612 20804 24668
rect 6626 24556 6636 24612
rect 6692 24556 11900 24612
rect 11956 24556 11966 24612
rect 14354 24556 14364 24612
rect 14420 24556 14980 24612
rect 15092 24556 16604 24612
rect 16660 24556 20804 24612
rect 21522 24556 21532 24612
rect 21588 24556 21868 24612
rect 21924 24556 21934 24612
rect 23314 24556 23324 24612
rect 23380 24556 23772 24612
rect 23828 24556 23838 24612
rect 26562 24556 26572 24612
rect 26628 24556 26908 24612
rect 26964 24556 26974 24612
rect 33954 24556 33964 24612
rect 34020 24556 34972 24612
rect 35028 24556 35038 24612
rect 36866 24556 36876 24612
rect 36932 24556 37996 24612
rect 38052 24556 40572 24612
rect 40628 24556 41692 24612
rect 41748 24556 41758 24612
rect 15092 24500 15148 24556
rect 1698 24444 1708 24500
rect 1764 24444 1774 24500
rect 10966 24444 11004 24500
rect 11060 24444 11070 24500
rect 12674 24444 12684 24500
rect 12740 24444 15148 24500
rect 18946 24444 18956 24500
rect 19012 24444 23212 24500
rect 23268 24444 23278 24500
rect 0 24276 800 24304
rect 1708 24276 1764 24444
rect 18722 24332 18732 24388
rect 18788 24332 21756 24388
rect 21812 24332 21822 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 42924 24276 42980 24780
rect 43474 24444 43484 24500
rect 43540 24444 46172 24500
rect 46228 24444 46238 24500
rect 0 24220 1764 24276
rect 12898 24220 12908 24276
rect 12964 24220 13356 24276
rect 13412 24220 14924 24276
rect 14980 24220 14990 24276
rect 15922 24220 15932 24276
rect 15988 24220 17612 24276
rect 17668 24220 18396 24276
rect 18452 24220 18462 24276
rect 42924 24220 43148 24276
rect 43204 24220 43214 24276
rect 0 24192 800 24220
rect 43484 24164 43540 24444
rect 13906 24108 13916 24164
rect 13972 24108 17388 24164
rect 17444 24108 17454 24164
rect 17826 24108 17836 24164
rect 17892 24108 19628 24164
rect 19684 24108 22092 24164
rect 22148 24108 23772 24164
rect 23828 24108 23838 24164
rect 43026 24108 43036 24164
rect 43092 24108 43540 24164
rect 16034 23996 16044 24052
rect 16100 23996 18172 24052
rect 18228 23996 18508 24052
rect 18564 23996 18574 24052
rect 20738 23996 20748 24052
rect 20804 23996 21532 24052
rect 21588 23996 21598 24052
rect 31154 23996 31164 24052
rect 31220 23996 31948 24052
rect 31892 23940 31948 23996
rect 7298 23884 7308 23940
rect 7364 23884 8204 23940
rect 8260 23884 8270 23940
rect 15698 23884 15708 23940
rect 15764 23884 23996 23940
rect 24052 23884 24062 23940
rect 31892 23884 33404 23940
rect 33460 23884 33470 23940
rect 33730 23884 33740 23940
rect 33796 23884 36092 23940
rect 36148 23884 42252 23940
rect 42308 23884 42318 23940
rect 50082 23884 50092 23940
rect 50148 23884 55580 23940
rect 55636 23884 55646 23940
rect 9986 23772 9996 23828
rect 10052 23772 10062 23828
rect 11778 23772 11788 23828
rect 11844 23772 14196 23828
rect 14690 23772 14700 23828
rect 14756 23772 16828 23828
rect 16884 23772 16894 23828
rect 17378 23772 17388 23828
rect 17444 23772 19404 23828
rect 19460 23772 19470 23828
rect 20402 23772 20412 23828
rect 20468 23772 31612 23828
rect 31668 23772 31678 23828
rect 41122 23772 41132 23828
rect 41188 23772 42140 23828
rect 42196 23772 42206 23828
rect 9996 23604 10052 23772
rect 14140 23716 14196 23772
rect 11218 23660 11228 23716
rect 11284 23660 13916 23716
rect 13972 23660 13982 23716
rect 14140 23660 16828 23716
rect 16884 23660 16940 23716
rect 16996 23660 17006 23716
rect 21298 23660 21308 23716
rect 21364 23660 22428 23716
rect 22484 23660 22494 23716
rect 25442 23660 25452 23716
rect 25508 23660 31948 23716
rect 32004 23660 32014 23716
rect 35746 23660 35756 23716
rect 35812 23660 36988 23716
rect 37044 23660 37054 23716
rect 40236 23660 41804 23716
rect 41860 23660 41870 23716
rect 42466 23660 42476 23716
rect 42532 23660 45500 23716
rect 45556 23660 45566 23716
rect 40236 23604 40292 23660
rect 59200 23604 60000 23632
rect 9996 23548 17332 23604
rect 21858 23548 21868 23604
rect 21924 23548 31388 23604
rect 31444 23548 31454 23604
rect 31602 23548 31612 23604
rect 31668 23548 40292 23604
rect 41682 23548 41692 23604
rect 41748 23548 42364 23604
rect 42420 23548 42430 23604
rect 42690 23548 42700 23604
rect 42756 23548 45948 23604
rect 46004 23548 47292 23604
rect 47348 23548 47358 23604
rect 57922 23548 57932 23604
rect 57988 23548 60000 23604
rect 16258 23436 16268 23492
rect 16324 23436 16940 23492
rect 16996 23436 17006 23492
rect 17276 23380 17332 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 59200 23520 60000 23548
rect 22978 23436 22988 23492
rect 23044 23436 23436 23492
rect 23492 23436 23502 23492
rect 24434 23436 24444 23492
rect 24500 23436 25564 23492
rect 25620 23436 25630 23492
rect 10994 23324 11004 23380
rect 11060 23324 11676 23380
rect 11732 23324 11742 23380
rect 13906 23324 13916 23380
rect 13972 23324 14252 23380
rect 14308 23324 14318 23380
rect 17266 23324 17276 23380
rect 17332 23324 17342 23380
rect 17602 23324 17612 23380
rect 17668 23324 22428 23380
rect 22484 23324 22494 23380
rect 26422 23324 26460 23380
rect 26516 23324 26526 23380
rect 37202 23324 37212 23380
rect 37268 23324 38444 23380
rect 38500 23324 40908 23380
rect 40964 23324 40974 23380
rect 11330 23212 11340 23268
rect 11396 23212 26684 23268
rect 26740 23212 26750 23268
rect 27458 23212 27468 23268
rect 27524 23212 28364 23268
rect 28420 23212 29484 23268
rect 29540 23212 29550 23268
rect 44258 23212 44268 23268
rect 44324 23212 44940 23268
rect 44996 23212 46172 23268
rect 46228 23212 46238 23268
rect 9314 23100 9324 23156
rect 9380 23100 11004 23156
rect 11060 23100 11070 23156
rect 15092 23100 16268 23156
rect 16324 23100 16492 23156
rect 16548 23100 16558 23156
rect 16706 23100 16716 23156
rect 16772 23100 18060 23156
rect 18116 23100 18126 23156
rect 20290 23100 20300 23156
rect 20356 23100 21420 23156
rect 21476 23100 21486 23156
rect 24658 23100 24668 23156
rect 24724 23100 25676 23156
rect 25732 23100 27580 23156
rect 27636 23100 28140 23156
rect 28196 23100 28206 23156
rect 31266 23100 31276 23156
rect 31332 23100 32060 23156
rect 32116 23100 32126 23156
rect 32498 23100 32508 23156
rect 32564 23100 33628 23156
rect 33684 23100 34860 23156
rect 34916 23100 35196 23156
rect 35252 23100 35262 23156
rect 35970 23100 35980 23156
rect 36036 23100 38892 23156
rect 38948 23100 38958 23156
rect 47842 23100 47852 23156
rect 47908 23100 48748 23156
rect 48804 23100 49084 23156
rect 49140 23100 49150 23156
rect 15092 22932 15148 23100
rect 15586 22988 15596 23044
rect 15652 22988 16156 23044
rect 16212 22988 17052 23044
rect 17108 22988 17118 23044
rect 22754 22988 22764 23044
rect 22820 22988 25340 23044
rect 25396 22988 25406 23044
rect 33506 22988 33516 23044
rect 33572 22988 34300 23044
rect 34356 22988 38332 23044
rect 38388 22988 39116 23044
rect 39172 22988 39182 23044
rect 42914 22988 42924 23044
rect 42980 22988 44604 23044
rect 44660 22988 45388 23044
rect 45444 22988 45454 23044
rect 46834 22988 46844 23044
rect 46900 22988 48860 23044
rect 48916 22988 48926 23044
rect 5618 22876 5628 22932
rect 5684 22876 7196 22932
rect 7252 22876 10108 22932
rect 10164 22876 11564 22932
rect 11620 22876 15148 22932
rect 17266 22876 17276 22932
rect 17332 22876 19348 22932
rect 19292 22820 19348 22876
rect 11442 22764 11452 22820
rect 11508 22764 18172 22820
rect 18228 22764 18238 22820
rect 19282 22764 19292 22820
rect 19348 22764 20188 22820
rect 20244 22764 20254 22820
rect 26002 22764 26012 22820
rect 26068 22764 26572 22820
rect 26628 22764 26638 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 17042 22652 17052 22708
rect 17108 22652 23324 22708
rect 23380 22652 23390 22708
rect 23548 22652 26908 22708
rect 26964 22652 26974 22708
rect 23548 22596 23604 22652
rect 13794 22540 13804 22596
rect 13860 22540 18508 22596
rect 18564 22540 20972 22596
rect 21028 22540 21038 22596
rect 22978 22540 22988 22596
rect 23044 22540 23604 22596
rect 26562 22540 26572 22596
rect 26628 22540 29932 22596
rect 29988 22540 29998 22596
rect 9874 22428 9884 22484
rect 9940 22428 12236 22484
rect 12292 22428 12302 22484
rect 15810 22428 15820 22484
rect 15876 22428 16716 22484
rect 16772 22428 16782 22484
rect 17826 22428 17836 22484
rect 17892 22428 20748 22484
rect 20804 22428 20814 22484
rect 21186 22428 21196 22484
rect 21252 22428 31500 22484
rect 31556 22428 32396 22484
rect 32452 22428 33516 22484
rect 33572 22428 33582 22484
rect 36194 22428 36204 22484
rect 36260 22428 36270 22484
rect 37762 22428 37772 22484
rect 37828 22428 45276 22484
rect 45332 22428 45342 22484
rect 20748 22372 20804 22428
rect 36204 22372 36260 22428
rect 6066 22316 6076 22372
rect 6132 22316 6972 22372
rect 7028 22316 7038 22372
rect 7410 22316 7420 22372
rect 7476 22316 8540 22372
rect 8596 22316 8988 22372
rect 9044 22316 9054 22372
rect 11666 22316 11676 22372
rect 11732 22316 12460 22372
rect 12516 22316 12526 22372
rect 19170 22316 19180 22372
rect 19236 22316 19740 22372
rect 19796 22316 19806 22372
rect 20178 22316 20188 22372
rect 20244 22316 20412 22372
rect 20468 22316 20478 22372
rect 20748 22316 21420 22372
rect 21476 22316 22316 22372
rect 22372 22316 22382 22372
rect 23398 22316 23436 22372
rect 23492 22316 26460 22372
rect 26516 22316 26526 22372
rect 26674 22316 26684 22372
rect 26740 22316 27020 22372
rect 27076 22316 27086 22372
rect 34514 22316 34524 22372
rect 34580 22316 35980 22372
rect 36036 22316 36046 22372
rect 36204 22316 44940 22372
rect 44996 22316 45724 22372
rect 45780 22316 45790 22372
rect 51090 22316 51100 22372
rect 51156 22316 55580 22372
rect 55636 22316 55646 22372
rect 26460 22260 26516 22316
rect 13878 22204 13916 22260
rect 13972 22204 13982 22260
rect 15092 22204 16380 22260
rect 16436 22204 16446 22260
rect 18946 22204 18956 22260
rect 19012 22204 22988 22260
rect 23044 22204 23054 22260
rect 26460 22204 29260 22260
rect 29316 22204 29326 22260
rect 15092 22148 15148 22204
rect 35980 22148 36036 22316
rect 59200 22260 60000 22288
rect 36194 22204 36204 22260
rect 36260 22204 37436 22260
rect 37492 22204 37502 22260
rect 41906 22204 41916 22260
rect 41972 22204 41982 22260
rect 45042 22204 45052 22260
rect 45108 22204 46172 22260
rect 46228 22204 46238 22260
rect 58146 22204 58156 22260
rect 58212 22204 60000 22260
rect 6738 22092 6748 22148
rect 6804 22092 7532 22148
rect 7588 22092 15148 22148
rect 15698 22092 15708 22148
rect 15764 22092 20188 22148
rect 20244 22092 21644 22148
rect 21700 22092 21710 22148
rect 24882 22092 24892 22148
rect 24948 22092 26908 22148
rect 35980 22092 40796 22148
rect 40852 22092 40862 22148
rect 11330 21980 11340 22036
rect 11396 21980 11676 22036
rect 11732 21980 11742 22036
rect 18610 21980 18620 22036
rect 18676 21980 19628 22036
rect 19684 21980 19694 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 6514 21868 6524 21924
rect 6580 21868 6590 21924
rect 11554 21868 11564 21924
rect 11620 21868 12348 21924
rect 12404 21868 13468 21924
rect 13524 21868 13534 21924
rect 16594 21868 16604 21924
rect 16660 21868 17836 21924
rect 17892 21868 17902 21924
rect 20188 21868 25900 21924
rect 25956 21868 25966 21924
rect 26852 21868 26908 22092
rect 41916 22036 41972 22204
rect 59200 22176 60000 22204
rect 38546 21980 38556 22036
rect 38612 21980 41972 22036
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 26964 21868 26974 21924
rect 33842 21868 33852 21924
rect 33908 21868 37324 21924
rect 37380 21868 37390 21924
rect 6524 21812 6580 21868
rect 20188 21812 20244 21868
rect 6524 21756 11228 21812
rect 11284 21756 17724 21812
rect 17780 21756 17790 21812
rect 19954 21756 19964 21812
rect 20020 21756 20244 21812
rect 24322 21756 24332 21812
rect 24388 21756 26012 21812
rect 26068 21756 26078 21812
rect 26450 21756 26460 21812
rect 26516 21756 31164 21812
rect 31220 21756 31230 21812
rect 31378 21756 31388 21812
rect 31444 21756 31948 21812
rect 32162 21756 32172 21812
rect 32228 21756 34972 21812
rect 35028 21756 35038 21812
rect 42466 21756 42476 21812
rect 42532 21756 43036 21812
rect 43092 21756 43102 21812
rect 31892 21700 31948 21756
rect 6514 21644 6524 21700
rect 6580 21644 8428 21700
rect 8484 21644 8494 21700
rect 11554 21644 11564 21700
rect 11620 21644 14140 21700
rect 14196 21644 14206 21700
rect 14354 21644 14364 21700
rect 14420 21644 20356 21700
rect 21074 21644 21084 21700
rect 21140 21644 23548 21700
rect 23604 21644 23614 21700
rect 26002 21644 26012 21700
rect 26068 21644 26236 21700
rect 26292 21644 26302 21700
rect 29810 21644 29820 21700
rect 29876 21644 31052 21700
rect 31108 21644 31118 21700
rect 31892 21644 43372 21700
rect 43428 21644 43438 21700
rect 20300 21588 20356 21644
rect 41580 21588 41636 21644
rect 59200 21588 60000 21616
rect 6626 21532 6636 21588
rect 6692 21532 7308 21588
rect 7364 21532 8092 21588
rect 8148 21532 8158 21588
rect 13122 21532 13132 21588
rect 13188 21532 13692 21588
rect 13748 21532 16156 21588
rect 16212 21532 16222 21588
rect 18610 21532 18620 21588
rect 18676 21532 18844 21588
rect 18900 21532 18910 21588
rect 20290 21532 20300 21588
rect 20356 21532 20366 21588
rect 22418 21532 22428 21588
rect 22484 21532 23100 21588
rect 23156 21532 23166 21588
rect 23426 21532 23436 21588
rect 23492 21532 25340 21588
rect 25396 21532 25406 21588
rect 33842 21532 33852 21588
rect 33908 21532 35084 21588
rect 35140 21532 35644 21588
rect 35700 21532 35710 21588
rect 36306 21532 36316 21588
rect 36372 21532 38556 21588
rect 38612 21532 38622 21588
rect 41570 21532 41580 21588
rect 41636 21532 41646 21588
rect 57922 21532 57932 21588
rect 57988 21532 60000 21588
rect 36316 21476 36372 21532
rect 59200 21504 60000 21532
rect 7858 21420 7868 21476
rect 7924 21420 8988 21476
rect 9044 21420 9054 21476
rect 10882 21420 10892 21476
rect 10948 21420 13356 21476
rect 13412 21420 15148 21476
rect 18274 21420 18284 21476
rect 18340 21420 19068 21476
rect 19124 21420 19134 21476
rect 19282 21420 19292 21476
rect 19348 21420 21868 21476
rect 21924 21420 21934 21476
rect 23846 21420 23884 21476
rect 23940 21420 23950 21476
rect 26786 21420 26796 21476
rect 26852 21420 27244 21476
rect 27300 21420 27310 21476
rect 29138 21420 29148 21476
rect 29204 21420 30604 21476
rect 30660 21420 30670 21476
rect 34626 21420 34636 21476
rect 34692 21420 36372 21476
rect 15092 21364 15148 21420
rect 15092 21308 15372 21364
rect 15428 21308 15438 21364
rect 18834 21308 18844 21364
rect 18900 21308 21532 21364
rect 21588 21308 21598 21364
rect 24210 21308 24220 21364
rect 24276 21308 31948 21364
rect 32498 21308 32508 21364
rect 32564 21308 35084 21364
rect 35140 21308 35150 21364
rect 31892 21252 31948 21308
rect 7858 21196 7868 21252
rect 7924 21196 11788 21252
rect 11844 21196 12572 21252
rect 12628 21196 12638 21252
rect 18946 21196 18956 21252
rect 19012 21196 19964 21252
rect 20020 21196 20030 21252
rect 31154 21196 31164 21252
rect 31220 21196 31612 21252
rect 31668 21196 31678 21252
rect 31892 21196 33516 21252
rect 33572 21196 33582 21252
rect 39330 21196 39340 21252
rect 39396 21196 41132 21252
rect 41188 21196 41198 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 9762 21084 9772 21140
rect 9828 21084 12236 21140
rect 12292 21084 12684 21140
rect 12740 21084 12750 21140
rect 18162 21084 18172 21140
rect 18228 21084 21084 21140
rect 21140 21084 21150 21140
rect 26226 21084 26236 21140
rect 26292 21084 26684 21140
rect 26740 21084 26750 21140
rect 12002 20972 12012 21028
rect 12068 20972 15148 21028
rect 15204 20972 15214 21028
rect 16706 20972 16716 21028
rect 16772 20972 25228 21028
rect 25284 20972 25294 21028
rect 32386 20972 32396 21028
rect 32452 20972 38108 21028
rect 38164 20972 38668 21028
rect 38724 20972 38734 21028
rect 0 20916 800 20944
rect 0 20860 1708 20916
rect 1764 20860 1774 20916
rect 14578 20860 14588 20916
rect 14644 20860 15036 20916
rect 15092 20860 17668 20916
rect 25666 20860 25676 20916
rect 25732 20860 29148 20916
rect 29204 20860 29214 20916
rect 34738 20860 34748 20916
rect 34804 20860 35868 20916
rect 35924 20860 35934 20916
rect 41346 20860 41356 20916
rect 41412 20860 42364 20916
rect 42420 20860 43148 20916
rect 43204 20860 43214 20916
rect 44034 20860 44044 20916
rect 44100 20860 47292 20916
rect 47348 20860 47358 20916
rect 48626 20860 48636 20916
rect 48692 20860 49532 20916
rect 49588 20860 49598 20916
rect 0 20832 800 20860
rect 17612 20804 17668 20860
rect 8306 20748 8316 20804
rect 8372 20748 9324 20804
rect 9380 20748 10220 20804
rect 10276 20748 10780 20804
rect 10836 20748 11788 20804
rect 11844 20748 11854 20804
rect 15092 20748 15372 20804
rect 15428 20748 15438 20804
rect 17602 20748 17612 20804
rect 17668 20748 17678 20804
rect 17938 20748 17948 20804
rect 18004 20748 18732 20804
rect 18788 20748 19404 20804
rect 19460 20748 19470 20804
rect 20598 20748 20636 20804
rect 20692 20748 20702 20804
rect 25330 20748 25340 20804
rect 25396 20748 28476 20804
rect 28532 20748 29820 20804
rect 29876 20748 29886 20804
rect 30930 20748 30940 20804
rect 30996 20748 31948 20804
rect 32004 20748 32284 20804
rect 32340 20748 32350 20804
rect 40226 20748 40236 20804
rect 40292 20748 41580 20804
rect 41636 20748 42756 20804
rect 46946 20748 46956 20804
rect 47012 20748 47964 20804
rect 48020 20748 48030 20804
rect 6290 20636 6300 20692
rect 6356 20636 10108 20692
rect 10164 20636 10174 20692
rect 12226 20636 12236 20692
rect 12292 20636 13468 20692
rect 13524 20636 14140 20692
rect 14196 20636 14206 20692
rect 15092 20580 15148 20748
rect 16594 20636 16604 20692
rect 16660 20636 26012 20692
rect 26068 20636 26078 20692
rect 27234 20636 27244 20692
rect 27300 20636 27692 20692
rect 27748 20636 31052 20692
rect 31108 20636 31118 20692
rect 31938 20636 31948 20692
rect 32004 20636 41468 20692
rect 41524 20636 41534 20692
rect 42700 20580 42756 20748
rect 46162 20636 46172 20692
rect 46228 20636 48860 20692
rect 48916 20636 48926 20692
rect 8642 20524 8652 20580
rect 8708 20524 13692 20580
rect 13748 20524 15148 20580
rect 16706 20524 16716 20580
rect 16772 20524 19852 20580
rect 19908 20524 20412 20580
rect 20468 20524 20478 20580
rect 20626 20524 20636 20580
rect 20692 20524 22540 20580
rect 22596 20524 22606 20580
rect 24518 20524 24556 20580
rect 24612 20524 24622 20580
rect 25228 20524 33852 20580
rect 33908 20524 33918 20580
rect 41122 20524 41132 20580
rect 41188 20524 41580 20580
rect 41636 20524 41646 20580
rect 42690 20524 42700 20580
rect 42756 20524 42766 20580
rect 9202 20412 9212 20468
rect 9268 20412 15148 20468
rect 17714 20412 17724 20468
rect 17780 20412 18844 20468
rect 18900 20412 18910 20468
rect 19282 20412 19292 20468
rect 19348 20412 19404 20468
rect 19460 20412 19470 20468
rect 21634 20412 21644 20468
rect 21700 20412 22764 20468
rect 22820 20412 25004 20468
rect 25060 20412 25070 20468
rect 15092 20356 15148 20412
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 25228 20356 25284 20524
rect 26786 20412 26796 20468
rect 26852 20412 31948 20468
rect 32004 20412 32014 20468
rect 32162 20412 32172 20468
rect 32228 20412 33516 20468
rect 33572 20412 33582 20468
rect 44034 20412 44044 20468
rect 44100 20412 45612 20468
rect 45668 20412 45678 20468
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 11862 20300 11900 20356
rect 11956 20300 11966 20356
rect 15092 20300 16268 20356
rect 16324 20300 17388 20356
rect 17444 20300 17454 20356
rect 17826 20300 17836 20356
rect 17892 20300 19460 20356
rect 22418 20300 22428 20356
rect 22484 20300 25284 20356
rect 27570 20300 27580 20356
rect 27636 20300 28364 20356
rect 28420 20300 28430 20356
rect 30716 20300 34748 20356
rect 34804 20300 34814 20356
rect 40898 20300 40908 20356
rect 40964 20300 43988 20356
rect 19404 20244 19460 20300
rect 30716 20244 30772 20300
rect 43932 20244 43988 20300
rect 6962 20188 6972 20244
rect 7028 20188 7038 20244
rect 7970 20188 7980 20244
rect 8036 20188 12068 20244
rect 12646 20188 12684 20244
rect 12740 20188 19180 20244
rect 19236 20188 19246 20244
rect 19404 20188 25340 20244
rect 25396 20188 25406 20244
rect 30706 20188 30716 20244
rect 30772 20188 30782 20244
rect 31714 20188 31724 20244
rect 31780 20188 33292 20244
rect 33348 20188 33358 20244
rect 41906 20188 41916 20244
rect 41972 20188 43708 20244
rect 43764 20188 43774 20244
rect 43922 20188 43932 20244
rect 43988 20188 44940 20244
rect 44996 20188 45006 20244
rect 58146 20188 58156 20244
rect 58212 20188 59332 20244
rect 6972 20132 7028 20188
rect 12012 20132 12068 20188
rect 6972 20076 7308 20132
rect 7364 20076 9156 20132
rect 11554 20076 11564 20132
rect 11620 20076 11676 20132
rect 11732 20076 11742 20132
rect 12002 20076 12012 20132
rect 12068 20076 12078 20132
rect 12572 20076 14812 20132
rect 14868 20076 14878 20132
rect 15138 20076 15148 20132
rect 15204 20076 15372 20132
rect 15428 20076 15438 20132
rect 15810 20076 15820 20132
rect 15876 20076 18060 20132
rect 18116 20076 18126 20132
rect 20402 20076 20412 20132
rect 20468 20076 22428 20132
rect 22484 20076 22494 20132
rect 24210 20076 24220 20132
rect 24276 20076 26236 20132
rect 26292 20076 26302 20132
rect 26852 20076 27468 20132
rect 27524 20076 27534 20132
rect 28130 20076 28140 20132
rect 28196 20076 28588 20132
rect 28644 20076 28654 20132
rect 33618 20076 33628 20132
rect 33684 20076 34076 20132
rect 34132 20076 34142 20132
rect 34962 20076 34972 20132
rect 35028 20076 37884 20132
rect 37940 20076 40124 20132
rect 40180 20076 40190 20132
rect 45938 20076 45948 20132
rect 46004 20076 47068 20132
rect 47124 20076 49196 20132
rect 49252 20076 49262 20132
rect 9100 20020 9156 20076
rect 12572 20020 12628 20076
rect 26852 20020 26908 20076
rect 5842 19964 5852 20020
rect 5908 19964 7084 20020
rect 7140 19964 7532 20020
rect 7588 19964 7598 20020
rect 8082 19964 8092 20020
rect 8148 19964 8540 20020
rect 8596 19964 8606 20020
rect 9100 19964 11452 20020
rect 11508 19964 12628 20020
rect 12898 19964 12908 20020
rect 12964 19964 13692 20020
rect 13748 19964 13758 20020
rect 14466 19964 14476 20020
rect 14532 19964 16716 20020
rect 16772 19964 16782 20020
rect 16930 19964 16940 20020
rect 16996 19964 17612 20020
rect 17668 19964 18620 20020
rect 18676 19964 18686 20020
rect 23426 19964 23436 20020
rect 23492 19964 25228 20020
rect 25284 19964 26908 20020
rect 27468 20020 27524 20076
rect 27468 19964 30044 20020
rect 30100 19964 30110 20020
rect 34514 19964 34524 20020
rect 34580 19964 36540 20020
rect 36596 19964 36606 20020
rect 39330 19964 39340 20020
rect 39396 19964 40460 20020
rect 40516 19964 40526 20020
rect 41682 19964 41692 20020
rect 41748 19964 42924 20020
rect 42980 19964 42990 20020
rect 11330 19852 11340 19908
rect 11396 19852 11676 19908
rect 11732 19852 12796 19908
rect 12852 19852 12862 19908
rect 15586 19852 15596 19908
rect 15652 19852 17500 19908
rect 17556 19852 20860 19908
rect 20916 19852 20926 19908
rect 26002 19852 26012 19908
rect 26068 19852 26908 19908
rect 27570 19852 27580 19908
rect 27636 19852 28924 19908
rect 28980 19852 28990 19908
rect 34290 19852 34300 19908
rect 34356 19852 37436 19908
rect 37492 19852 37502 19908
rect 40002 19852 40012 19908
rect 40068 19852 43596 19908
rect 43652 19852 45948 19908
rect 46004 19852 46014 19908
rect 26852 19796 26908 19852
rect 59276 19796 59332 20188
rect 8754 19740 8764 19796
rect 8820 19740 12572 19796
rect 12628 19740 12638 19796
rect 13906 19740 13916 19796
rect 13972 19740 17500 19796
rect 17556 19740 17566 19796
rect 18162 19740 18172 19796
rect 18228 19740 19292 19796
rect 19348 19740 20076 19796
rect 20132 19740 21420 19796
rect 21476 19740 25452 19796
rect 25508 19740 25518 19796
rect 25778 19740 25788 19796
rect 25844 19740 26236 19796
rect 26292 19740 26302 19796
rect 26852 19740 33628 19796
rect 33684 19740 33694 19796
rect 35970 19740 35980 19796
rect 36036 19740 37660 19796
rect 37716 19740 38332 19796
rect 38388 19740 38398 19796
rect 43698 19740 43708 19796
rect 43764 19740 46284 19796
rect 46340 19740 47964 19796
rect 48020 19740 48972 19796
rect 49028 19740 49308 19796
rect 49364 19740 49374 19796
rect 59052 19740 59332 19796
rect 9996 19628 14364 19684
rect 14420 19628 14430 19684
rect 16594 19628 16604 19684
rect 16660 19628 26740 19684
rect 31938 19628 31948 19684
rect 32004 19628 33740 19684
rect 33796 19628 33806 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 7074 19292 7084 19348
rect 7140 19292 7756 19348
rect 7812 19292 7822 19348
rect 9996 19236 10052 19628
rect 26684 19572 26740 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 59052 19572 59108 19740
rect 59200 19572 60000 19600
rect 13458 19516 13468 19572
rect 13524 19516 23996 19572
rect 24052 19516 24062 19572
rect 24210 19516 24220 19572
rect 24276 19516 25676 19572
rect 25732 19516 26460 19572
rect 26516 19516 26526 19572
rect 26674 19516 26684 19572
rect 26740 19516 28140 19572
rect 28196 19516 29148 19572
rect 29204 19516 29932 19572
rect 29988 19516 30380 19572
rect 30436 19516 30446 19572
rect 59052 19516 60000 19572
rect 59200 19488 60000 19516
rect 10630 19404 10668 19460
rect 10724 19404 10734 19460
rect 10994 19404 11004 19460
rect 11060 19404 16604 19460
rect 16660 19404 16670 19460
rect 17154 19404 17164 19460
rect 17220 19404 18172 19460
rect 18228 19404 18238 19460
rect 18386 19404 18396 19460
rect 18452 19404 22988 19460
rect 23044 19404 23054 19460
rect 40674 19404 40684 19460
rect 40740 19404 41692 19460
rect 41748 19404 41758 19460
rect 10210 19292 10220 19348
rect 10276 19292 14476 19348
rect 14532 19292 14542 19348
rect 15026 19292 15036 19348
rect 15092 19292 21980 19348
rect 22036 19292 22316 19348
rect 22372 19292 22382 19348
rect 25106 19292 25116 19348
rect 25172 19292 27132 19348
rect 27188 19292 27198 19348
rect 31266 19292 31276 19348
rect 31332 19292 31612 19348
rect 31668 19292 32732 19348
rect 32788 19292 33068 19348
rect 33124 19292 33134 19348
rect 38546 19292 38556 19348
rect 38612 19292 38622 19348
rect 38556 19236 38612 19292
rect 6738 19180 6748 19236
rect 6804 19180 7308 19236
rect 7364 19180 7374 19236
rect 9090 19180 9100 19236
rect 9156 19180 9324 19236
rect 9380 19180 9390 19236
rect 9650 19180 9660 19236
rect 9716 19180 10052 19236
rect 12002 19180 12012 19236
rect 12068 19180 14252 19236
rect 14308 19180 14812 19236
rect 14868 19180 14878 19236
rect 18722 19180 18732 19236
rect 18788 19180 19068 19236
rect 19124 19180 19292 19236
rect 19348 19180 19358 19236
rect 20402 19180 20412 19236
rect 20468 19180 22876 19236
rect 22932 19180 22942 19236
rect 25974 19180 26012 19236
rect 26068 19180 26078 19236
rect 26226 19180 26236 19236
rect 26292 19180 28476 19236
rect 28532 19180 28542 19236
rect 30930 19180 30940 19236
rect 30996 19180 38332 19236
rect 38388 19180 38612 19236
rect 50418 19180 50428 19236
rect 50484 19180 51436 19236
rect 51492 19180 51502 19236
rect 7074 19068 7084 19124
rect 7140 19068 9884 19124
rect 9940 19068 9950 19124
rect 10882 19068 10892 19124
rect 10948 19068 12236 19124
rect 12292 19068 12302 19124
rect 14018 19068 14028 19124
rect 14084 19068 15036 19124
rect 15092 19068 15708 19124
rect 15764 19068 15774 19124
rect 16380 19068 17052 19124
rect 17108 19068 17164 19124
rect 17220 19068 17230 19124
rect 17490 19068 17500 19124
rect 17556 19068 20916 19124
rect 22306 19068 22316 19124
rect 22372 19068 22652 19124
rect 22708 19068 22718 19124
rect 23538 19068 23548 19124
rect 23604 19068 23884 19124
rect 23940 19068 23950 19124
rect 49522 19068 49532 19124
rect 49588 19068 50204 19124
rect 50260 19068 50270 19124
rect 16380 19012 16436 19068
rect 20860 19012 20916 19068
rect 8642 18956 8652 19012
rect 8708 18956 9548 19012
rect 9604 18956 9614 19012
rect 12562 18956 12572 19012
rect 12628 18956 16436 19012
rect 16594 18956 16604 19012
rect 16660 18956 18620 19012
rect 18676 18956 19180 19012
rect 19236 18956 19246 19012
rect 20402 18956 20412 19012
rect 20468 18956 20478 19012
rect 20860 18956 25228 19012
rect 25284 18956 25294 19012
rect 25442 18956 25452 19012
rect 25508 18956 31612 19012
rect 31668 18956 31678 19012
rect 33954 18956 33964 19012
rect 34020 18956 34524 19012
rect 34580 18956 34590 19012
rect 40786 18956 40796 19012
rect 40852 18956 41580 19012
rect 41636 18956 41646 19012
rect 8978 18844 8988 18900
rect 9044 18844 11676 18900
rect 11732 18844 13020 18900
rect 13076 18844 13086 18900
rect 13346 18844 13356 18900
rect 13412 18844 13748 18900
rect 13692 18676 13748 18844
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 20412 18788 20468 18956
rect 59200 18900 60000 18928
rect 22530 18844 22540 18900
rect 22596 18844 23324 18900
rect 23380 18844 27468 18900
rect 27524 18844 27534 18900
rect 36418 18844 36428 18900
rect 36484 18844 37212 18900
rect 37268 18844 39452 18900
rect 39508 18844 40124 18900
rect 40180 18844 40190 18900
rect 58146 18844 58156 18900
rect 58212 18844 60000 18900
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 59200 18816 60000 18844
rect 20412 18732 27132 18788
rect 27188 18732 28588 18788
rect 28644 18732 29260 18788
rect 29316 18732 29540 18788
rect 29484 18676 29540 18732
rect 5954 18620 5964 18676
rect 6020 18620 7756 18676
rect 7812 18620 7980 18676
rect 8036 18620 8046 18676
rect 8978 18620 8988 18676
rect 9044 18620 9436 18676
rect 9492 18620 9502 18676
rect 10546 18620 10556 18676
rect 10612 18620 11004 18676
rect 11060 18620 11070 18676
rect 11330 18620 11340 18676
rect 11396 18620 13468 18676
rect 13524 18620 13534 18676
rect 13692 18620 16828 18676
rect 16884 18620 16894 18676
rect 19394 18620 19404 18676
rect 19460 18620 21868 18676
rect 21924 18620 25004 18676
rect 25060 18620 25070 18676
rect 29474 18620 29484 18676
rect 29540 18620 29550 18676
rect 6514 18508 6524 18564
rect 6580 18508 8316 18564
rect 8372 18508 8382 18564
rect 8866 18508 8876 18564
rect 8932 18508 9772 18564
rect 9828 18508 10332 18564
rect 10388 18508 10398 18564
rect 11442 18508 11452 18564
rect 11508 18508 16100 18564
rect 16258 18508 16268 18564
rect 16324 18508 16380 18564
rect 16436 18508 16446 18564
rect 16678 18508 16716 18564
rect 16772 18508 16782 18564
rect 18834 18508 18844 18564
rect 18900 18508 23772 18564
rect 23828 18508 23838 18564
rect 27682 18508 27692 18564
rect 27748 18508 30492 18564
rect 30548 18508 30558 18564
rect 38546 18508 38556 18564
rect 38612 18508 44044 18564
rect 44100 18508 44716 18564
rect 44772 18508 44782 18564
rect 16044 18452 16100 18508
rect 6066 18396 6076 18452
rect 6132 18396 6748 18452
rect 6804 18396 6814 18452
rect 9314 18396 9324 18452
rect 9380 18396 10444 18452
rect 10500 18396 10510 18452
rect 13122 18396 13132 18452
rect 13188 18396 13692 18452
rect 13748 18396 13758 18452
rect 16044 18396 17388 18452
rect 17444 18396 17454 18452
rect 17602 18396 17612 18452
rect 17668 18396 18620 18452
rect 18676 18396 18686 18452
rect 19618 18396 19628 18452
rect 19684 18396 21308 18452
rect 21364 18396 21374 18452
rect 22418 18396 22428 18452
rect 22484 18396 22988 18452
rect 23044 18396 23436 18452
rect 23492 18396 23502 18452
rect 23772 18396 28812 18452
rect 28868 18396 28878 18452
rect 37090 18396 37100 18452
rect 37156 18396 37772 18452
rect 37828 18396 37838 18452
rect 38434 18396 38444 18452
rect 38500 18396 39228 18452
rect 39284 18396 39294 18452
rect 43250 18396 43260 18452
rect 43316 18396 46060 18452
rect 46116 18396 46126 18452
rect 48738 18396 48748 18452
rect 48804 18396 49644 18452
rect 49700 18396 49710 18452
rect 9762 18284 9772 18340
rect 9828 18284 10108 18340
rect 10164 18284 12684 18340
rect 12740 18284 12750 18340
rect 13570 18284 13580 18340
rect 13636 18284 17276 18340
rect 17332 18284 17342 18340
rect 17714 18284 17724 18340
rect 17780 18284 23324 18340
rect 23380 18284 23390 18340
rect 10434 18172 10444 18228
rect 10500 18172 10668 18228
rect 10724 18172 10734 18228
rect 10994 18172 11004 18228
rect 11060 18172 11340 18228
rect 11396 18172 11406 18228
rect 15250 18172 15260 18228
rect 15316 18172 19628 18228
rect 19684 18172 22540 18228
rect 22596 18172 22606 18228
rect 23324 18116 23380 18284
rect 23772 18228 23828 18396
rect 24546 18284 24556 18340
rect 24612 18284 25900 18340
rect 25956 18284 25966 18340
rect 27654 18284 27692 18340
rect 27748 18284 27758 18340
rect 38546 18284 38556 18340
rect 38612 18284 39340 18340
rect 39396 18284 39406 18340
rect 40114 18284 40124 18340
rect 40180 18284 45948 18340
rect 46004 18284 46014 18340
rect 50306 18284 50316 18340
rect 50372 18284 51660 18340
rect 51716 18284 51726 18340
rect 59200 18228 60000 18256
rect 23762 18172 23772 18228
rect 23828 18172 23838 18228
rect 25554 18172 25564 18228
rect 25620 18172 30604 18228
rect 30660 18172 30670 18228
rect 57922 18172 57932 18228
rect 57988 18172 60000 18228
rect 59200 18144 60000 18172
rect 9762 18060 9772 18116
rect 9828 18060 16604 18116
rect 16660 18060 16670 18116
rect 16930 18060 16940 18116
rect 16996 18060 19068 18116
rect 19124 18060 19134 18116
rect 19506 18060 19516 18116
rect 19572 18060 20188 18116
rect 20244 18060 20254 18116
rect 23324 18060 25004 18116
rect 25060 18060 25070 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 19068 18004 19124 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 6850 17948 6860 18004
rect 6916 17948 10052 18004
rect 10322 17948 10332 18004
rect 10388 17948 17612 18004
rect 17668 17948 17678 18004
rect 19068 17948 23772 18004
rect 23828 17948 23838 18004
rect 33394 17948 33404 18004
rect 33460 17948 34300 18004
rect 34356 17948 34366 18004
rect 9996 17892 10052 17948
rect 4386 17836 4396 17892
rect 4452 17836 8652 17892
rect 8708 17836 8718 17892
rect 9996 17836 15932 17892
rect 15988 17836 15998 17892
rect 18722 17836 18732 17892
rect 18788 17836 20412 17892
rect 20468 17836 20478 17892
rect 23286 17836 23324 17892
rect 23380 17836 23390 17892
rect 28242 17836 28252 17892
rect 28308 17836 34748 17892
rect 34804 17836 35756 17892
rect 35812 17836 36988 17892
rect 37044 17836 38444 17892
rect 38500 17836 38510 17892
rect 8652 17780 8708 17836
rect 7746 17724 7756 17780
rect 7812 17724 8092 17780
rect 8148 17724 8428 17780
rect 8484 17724 8494 17780
rect 8652 17724 11340 17780
rect 11396 17724 11676 17780
rect 11732 17724 11742 17780
rect 15810 17724 15820 17780
rect 15876 17724 19292 17780
rect 19348 17724 19628 17780
rect 19684 17724 19694 17780
rect 23762 17724 23772 17780
rect 23828 17724 25452 17780
rect 25508 17724 25518 17780
rect 25890 17724 25900 17780
rect 25956 17724 26236 17780
rect 26292 17724 26302 17780
rect 29698 17724 29708 17780
rect 29764 17724 32620 17780
rect 32676 17724 32686 17780
rect 35410 17724 35420 17780
rect 35476 17724 35980 17780
rect 36036 17724 36046 17780
rect 47506 17724 47516 17780
rect 47572 17724 49532 17780
rect 49588 17724 49598 17780
rect 5058 17612 5068 17668
rect 5124 17612 5740 17668
rect 5796 17612 5806 17668
rect 7298 17612 7308 17668
rect 7364 17612 8316 17668
rect 8372 17612 8382 17668
rect 10098 17612 10108 17668
rect 10164 17612 11004 17668
rect 11060 17612 16940 17668
rect 16996 17612 17006 17668
rect 17714 17612 17724 17668
rect 17780 17612 21980 17668
rect 22036 17612 22046 17668
rect 23538 17612 23548 17668
rect 23604 17612 24332 17668
rect 24388 17612 24398 17668
rect 26002 17612 26012 17668
rect 26068 17612 26908 17668
rect 26964 17612 26974 17668
rect 31892 17612 34300 17668
rect 34356 17612 35532 17668
rect 35588 17612 35598 17668
rect 41346 17612 41356 17668
rect 41412 17612 42700 17668
rect 42756 17612 42766 17668
rect 46498 17612 46508 17668
rect 46564 17612 47068 17668
rect 47124 17612 47134 17668
rect 47282 17612 47292 17668
rect 47348 17612 48076 17668
rect 48132 17612 48142 17668
rect 48626 17612 48636 17668
rect 48692 17612 49196 17668
rect 49252 17612 49262 17668
rect 50194 17612 50204 17668
rect 50260 17612 51324 17668
rect 51380 17612 51390 17668
rect 52994 17612 53004 17668
rect 53060 17612 55580 17668
rect 55636 17612 55646 17668
rect 0 17556 800 17584
rect 31892 17556 31948 17612
rect 48636 17556 48692 17612
rect 0 17500 1708 17556
rect 1764 17500 1774 17556
rect 9986 17500 9996 17556
rect 10052 17500 10668 17556
rect 10724 17500 10734 17556
rect 12898 17500 12908 17556
rect 12964 17500 15484 17556
rect 15540 17500 15550 17556
rect 17266 17500 17276 17556
rect 17332 17500 21420 17556
rect 21476 17500 21486 17556
rect 22978 17500 22988 17556
rect 23044 17500 26572 17556
rect 26628 17500 26638 17556
rect 31714 17500 31724 17556
rect 31780 17500 31948 17556
rect 33394 17500 33404 17556
rect 33460 17500 34076 17556
rect 34132 17500 34524 17556
rect 34580 17500 34590 17556
rect 43250 17500 43260 17556
rect 43316 17500 43708 17556
rect 46946 17500 46956 17556
rect 47012 17500 47404 17556
rect 47460 17500 48692 17556
rect 50082 17500 50092 17556
rect 50148 17500 50652 17556
rect 50708 17500 51100 17556
rect 51156 17500 51166 17556
rect 0 17472 800 17500
rect 43652 17444 43708 17500
rect 14438 17388 14476 17444
rect 14532 17388 14542 17444
rect 15092 17388 17724 17444
rect 17780 17388 17790 17444
rect 18610 17388 18620 17444
rect 18676 17388 24220 17444
rect 24276 17388 26908 17444
rect 26964 17388 26974 17444
rect 37202 17388 37212 17444
rect 37268 17388 38332 17444
rect 38388 17388 39116 17444
rect 39172 17388 40908 17444
rect 40964 17388 40974 17444
rect 43652 17388 44268 17444
rect 44324 17388 44334 17444
rect 15092 17332 15148 17388
rect 6962 17276 6972 17332
rect 7028 17276 9772 17332
rect 9828 17276 15148 17332
rect 16594 17276 16604 17332
rect 16660 17276 17388 17332
rect 17444 17276 17948 17332
rect 18004 17276 18014 17332
rect 20626 17276 20636 17332
rect 20692 17276 21532 17332
rect 21588 17276 21598 17332
rect 24546 17276 24556 17332
rect 24612 17276 27692 17332
rect 27748 17276 27758 17332
rect 41682 17276 41692 17332
rect 41748 17276 41916 17332
rect 41972 17276 41982 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 6066 17164 6076 17220
rect 6132 17164 13916 17220
rect 13972 17164 14476 17220
rect 14532 17164 14542 17220
rect 15922 17164 15932 17220
rect 15988 17164 17612 17220
rect 17668 17164 18508 17220
rect 18564 17164 18574 17220
rect 26226 17164 26236 17220
rect 26292 17164 27804 17220
rect 27860 17164 28364 17220
rect 28420 17164 28430 17220
rect 36978 17164 36988 17220
rect 37044 17164 37660 17220
rect 37716 17164 37726 17220
rect 5506 17052 5516 17108
rect 5572 17052 7084 17108
rect 7140 17052 7150 17108
rect 7410 17052 7420 17108
rect 7476 17052 7756 17108
rect 7812 17052 7822 17108
rect 11106 17052 11116 17108
rect 11172 17052 11564 17108
rect 11620 17052 11630 17108
rect 15138 17052 15148 17108
rect 15204 17052 15372 17108
rect 15428 17052 16156 17108
rect 16212 17052 16222 17108
rect 17938 17052 17948 17108
rect 18004 17052 23996 17108
rect 24052 17052 24332 17108
rect 24388 17052 24398 17108
rect 24546 17052 24556 17108
rect 24612 17052 27244 17108
rect 27300 17052 27310 17108
rect 41122 17052 41132 17108
rect 41188 17052 43372 17108
rect 43428 17052 43708 17108
rect 43652 16996 43708 17052
rect 6850 16940 6860 16996
rect 6916 16940 8428 16996
rect 8484 16940 8494 16996
rect 8642 16940 8652 16996
rect 8708 16940 10332 16996
rect 10388 16940 10398 16996
rect 14914 16940 14924 16996
rect 14980 16940 18172 16996
rect 18228 16940 18238 16996
rect 21186 16940 21196 16996
rect 21252 16940 23772 16996
rect 23828 16940 23838 16996
rect 24630 16940 24668 16996
rect 24724 16940 25788 16996
rect 25844 16940 25854 16996
rect 26226 16940 26236 16996
rect 26292 16940 28028 16996
rect 28084 16940 30492 16996
rect 30548 16940 31052 16996
rect 31108 16940 31118 16996
rect 36082 16940 36092 16996
rect 36148 16940 37660 16996
rect 37716 16940 37726 16996
rect 43652 16940 43820 16996
rect 43876 16940 44604 16996
rect 44660 16940 46844 16996
rect 46900 16940 46910 16996
rect 59200 16884 60000 16912
rect 6738 16828 6748 16884
rect 6804 16828 7756 16884
rect 7812 16828 7822 16884
rect 9986 16828 9996 16884
rect 10052 16828 13580 16884
rect 13636 16828 13916 16884
rect 13972 16828 13982 16884
rect 15362 16828 15372 16884
rect 15428 16828 15932 16884
rect 15988 16828 15998 16884
rect 16818 16828 16828 16884
rect 16884 16828 17948 16884
rect 18004 16828 18014 16884
rect 19740 16828 20860 16884
rect 20916 16828 20926 16884
rect 23090 16828 23100 16884
rect 23156 16828 27132 16884
rect 27188 16828 31164 16884
rect 31220 16828 31230 16884
rect 34402 16828 34412 16884
rect 34468 16828 36428 16884
rect 36484 16828 36494 16884
rect 36754 16828 36764 16884
rect 36820 16828 37212 16884
rect 37268 16828 37278 16884
rect 41010 16828 41020 16884
rect 41076 16828 41636 16884
rect 41794 16828 41804 16884
rect 41860 16828 42588 16884
rect 42644 16828 42654 16884
rect 43362 16828 43372 16884
rect 43428 16828 47516 16884
rect 47572 16828 47582 16884
rect 51874 16828 51884 16884
rect 51940 16828 53116 16884
rect 53172 16828 53182 16884
rect 58044 16828 60000 16884
rect 19740 16772 19796 16828
rect 41580 16772 41636 16828
rect 58044 16772 58100 16828
rect 59200 16800 60000 16828
rect 13458 16716 13468 16772
rect 13524 16716 19404 16772
rect 19460 16716 19470 16772
rect 19628 16716 19796 16772
rect 19852 16716 27468 16772
rect 27524 16716 29708 16772
rect 29764 16716 29774 16772
rect 41580 16716 41916 16772
rect 41972 16716 41982 16772
rect 57922 16716 57932 16772
rect 57988 16716 58100 16772
rect 19628 16660 19684 16716
rect 19852 16660 19908 16716
rect 11190 16604 11228 16660
rect 11284 16604 11294 16660
rect 11890 16604 11900 16660
rect 11956 16604 19684 16660
rect 19842 16604 19852 16660
rect 19908 16604 19918 16660
rect 26786 16604 26796 16660
rect 26852 16604 31836 16660
rect 31892 16604 31902 16660
rect 36306 16604 36316 16660
rect 36372 16604 40796 16660
rect 40852 16604 41468 16660
rect 41524 16604 41534 16660
rect 46834 16604 46844 16660
rect 46900 16604 47628 16660
rect 47684 16604 47694 16660
rect 13682 16492 13692 16548
rect 13748 16492 14924 16548
rect 14980 16492 14990 16548
rect 16818 16492 16828 16548
rect 16884 16492 17948 16548
rect 18004 16492 18014 16548
rect 19170 16492 19180 16548
rect 19236 16492 21868 16548
rect 21924 16492 21934 16548
rect 28690 16492 28700 16548
rect 28756 16492 29260 16548
rect 29316 16492 29326 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 4946 16380 4956 16436
rect 5012 16380 5516 16436
rect 5572 16380 7420 16436
rect 7476 16380 12348 16436
rect 12404 16380 12414 16436
rect 14578 16380 14588 16436
rect 14644 16380 15036 16436
rect 15092 16380 15102 16436
rect 17462 16380 17500 16436
rect 17556 16380 17566 16436
rect 20514 16380 20524 16436
rect 20580 16380 20636 16436
rect 20692 16380 20702 16436
rect 25106 16380 25116 16436
rect 25172 16380 31948 16436
rect 31892 16324 31948 16380
rect 6626 16268 6636 16324
rect 6692 16268 9660 16324
rect 9716 16268 9726 16324
rect 14914 16268 14924 16324
rect 14980 16268 18844 16324
rect 18900 16268 18910 16324
rect 19954 16268 19964 16324
rect 20020 16268 21644 16324
rect 21700 16268 21710 16324
rect 25330 16268 25340 16324
rect 25396 16268 26684 16324
rect 26740 16268 26796 16324
rect 26852 16268 26862 16324
rect 31892 16268 41356 16324
rect 41412 16268 41422 16324
rect 41906 16268 41916 16324
rect 41972 16268 45388 16324
rect 45444 16268 45454 16324
rect 59200 16212 60000 16240
rect 8866 16156 8876 16212
rect 8932 16156 9940 16212
rect 11330 16156 11340 16212
rect 11396 16156 13356 16212
rect 13412 16156 13422 16212
rect 15250 16156 15260 16212
rect 15316 16156 15484 16212
rect 15540 16156 16492 16212
rect 16548 16156 16558 16212
rect 17154 16156 17164 16212
rect 17220 16156 18060 16212
rect 18116 16156 19292 16212
rect 19348 16156 19358 16212
rect 19730 16156 19740 16212
rect 19796 16156 22316 16212
rect 22372 16156 22382 16212
rect 23426 16156 23436 16212
rect 23492 16156 25564 16212
rect 25620 16156 25630 16212
rect 27570 16156 27580 16212
rect 27636 16156 27916 16212
rect 27972 16156 27982 16212
rect 29698 16156 29708 16212
rect 29764 16156 30380 16212
rect 30436 16156 30446 16212
rect 33394 16156 33404 16212
rect 33460 16156 33964 16212
rect 34020 16156 34412 16212
rect 34468 16156 34478 16212
rect 35970 16156 35980 16212
rect 36036 16156 37436 16212
rect 37492 16156 37502 16212
rect 39228 16156 45724 16212
rect 45780 16156 45790 16212
rect 50194 16156 50204 16212
rect 50260 16156 51212 16212
rect 51268 16156 51278 16212
rect 58146 16156 58156 16212
rect 58212 16156 60000 16212
rect 9884 16100 9940 16156
rect 39228 16100 39284 16156
rect 59200 16128 60000 16156
rect 7522 16044 7532 16100
rect 7588 16044 9548 16100
rect 9604 16044 9614 16100
rect 9874 16044 9884 16100
rect 9940 16044 13580 16100
rect 13636 16044 13646 16100
rect 16930 16044 16940 16100
rect 16996 16044 22428 16100
rect 22484 16044 22494 16100
rect 22754 16044 22764 16100
rect 22820 16044 23324 16100
rect 23380 16044 23390 16100
rect 23874 16044 23884 16100
rect 23940 16044 25004 16100
rect 25060 16044 25070 16100
rect 26674 16044 26684 16100
rect 26740 16044 27804 16100
rect 27860 16044 27870 16100
rect 33506 16044 33516 16100
rect 33572 16044 34300 16100
rect 34356 16044 34366 16100
rect 35186 16044 35196 16100
rect 35252 16044 39284 16100
rect 40114 16044 40124 16100
rect 40180 16044 41356 16100
rect 41412 16044 41422 16100
rect 50082 16044 50092 16100
rect 50148 16044 50876 16100
rect 50932 16044 50942 16100
rect 52994 16044 53004 16100
rect 53060 16044 55580 16100
rect 55636 16044 55646 16100
rect 4722 15932 4732 15988
rect 4788 15932 9212 15988
rect 9268 15932 10444 15988
rect 10500 15932 10510 15988
rect 14466 15932 14476 15988
rect 14532 15932 21812 15988
rect 21970 15932 21980 15988
rect 22036 15932 28924 15988
rect 28980 15932 29484 15988
rect 29540 15932 29550 15988
rect 32946 15932 32956 15988
rect 33012 15932 33628 15988
rect 33684 15932 33694 15988
rect 34066 15932 34076 15988
rect 34132 15932 35756 15988
rect 35812 15932 35822 15988
rect 51538 15932 51548 15988
rect 51604 15932 52668 15988
rect 52724 15932 52734 15988
rect 21756 15876 21812 15932
rect 14018 15820 14028 15876
rect 14084 15820 16940 15876
rect 16996 15820 17006 15876
rect 17164 15820 17612 15876
rect 17668 15820 20524 15876
rect 20580 15820 20590 15876
rect 21756 15820 22092 15876
rect 22148 15820 22988 15876
rect 23044 15820 23054 15876
rect 23958 15820 23996 15876
rect 24052 15820 24062 15876
rect 24434 15820 24444 15876
rect 24500 15820 25116 15876
rect 25172 15820 25182 15876
rect 27122 15820 27132 15876
rect 27188 15820 29036 15876
rect 29092 15820 29102 15876
rect 29810 15820 29820 15876
rect 29876 15820 30828 15876
rect 30884 15820 30894 15876
rect 31714 15820 31724 15876
rect 31780 15820 33180 15876
rect 33236 15820 33246 15876
rect 38210 15820 38220 15876
rect 38276 15820 39900 15876
rect 39956 15820 39966 15876
rect 41458 15820 41468 15876
rect 41524 15820 42364 15876
rect 42420 15820 42430 15876
rect 49858 15820 49868 15876
rect 49924 15820 50988 15876
rect 51044 15820 51054 15876
rect 17164 15764 17220 15820
rect 8082 15708 8092 15764
rect 8148 15708 12572 15764
rect 12628 15708 12638 15764
rect 13570 15708 13580 15764
rect 13636 15708 17220 15764
rect 21942 15708 21980 15764
rect 22036 15708 22046 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 5954 15596 5964 15652
rect 6020 15596 14140 15652
rect 14196 15596 15036 15652
rect 15092 15596 15102 15652
rect 21410 15596 21420 15652
rect 21476 15596 22540 15652
rect 22596 15596 25788 15652
rect 25844 15596 25854 15652
rect 27682 15596 27692 15652
rect 27748 15596 28588 15652
rect 28644 15596 28654 15652
rect 31490 15596 31500 15652
rect 31556 15596 31612 15652
rect 31668 15596 31678 15652
rect 59200 15540 60000 15568
rect 5058 15484 5068 15540
rect 5124 15484 11452 15540
rect 11508 15484 11518 15540
rect 11778 15484 11788 15540
rect 11844 15484 11882 15540
rect 13122 15484 13132 15540
rect 13188 15484 14252 15540
rect 14308 15484 18172 15540
rect 18228 15484 19628 15540
rect 19684 15484 21308 15540
rect 21364 15484 21374 15540
rect 24434 15484 24444 15540
rect 24500 15484 24668 15540
rect 24724 15484 24734 15540
rect 28130 15484 28140 15540
rect 28196 15484 29372 15540
rect 29428 15484 29438 15540
rect 34066 15484 34076 15540
rect 34132 15484 35084 15540
rect 35140 15484 35150 15540
rect 57922 15484 57932 15540
rect 57988 15484 60000 15540
rect 59200 15456 60000 15484
rect 8754 15372 8764 15428
rect 8820 15372 9324 15428
rect 9380 15372 9390 15428
rect 10770 15372 10780 15428
rect 10836 15372 14924 15428
rect 14980 15372 14990 15428
rect 15082 15372 15092 15428
rect 15148 15372 15764 15428
rect 16930 15372 16940 15428
rect 16996 15372 17052 15428
rect 17108 15372 17118 15428
rect 17378 15372 17388 15428
rect 17444 15372 19124 15428
rect 19282 15372 19292 15428
rect 19348 15372 19740 15428
rect 19796 15372 19806 15428
rect 21382 15372 21420 15428
rect 21476 15372 21486 15428
rect 22754 15372 22764 15428
rect 22820 15372 22830 15428
rect 24658 15372 24668 15428
rect 24724 15372 26012 15428
rect 26068 15372 26078 15428
rect 26898 15372 26908 15428
rect 26964 15372 27580 15428
rect 27636 15372 27646 15428
rect 48290 15372 48300 15428
rect 48356 15372 51100 15428
rect 51156 15372 52332 15428
rect 52388 15372 52398 15428
rect 7298 15260 7308 15316
rect 7364 15260 13692 15316
rect 13748 15260 13758 15316
rect 14242 15260 14252 15316
rect 14308 15260 15484 15316
rect 15540 15260 15550 15316
rect 15708 15204 15764 15372
rect 19068 15316 19124 15372
rect 22764 15316 22820 15372
rect 17938 15260 17948 15316
rect 18004 15260 18732 15316
rect 18788 15260 18798 15316
rect 19068 15260 22764 15316
rect 22820 15260 22830 15316
rect 26562 15260 26572 15316
rect 26628 15260 26908 15316
rect 27906 15260 27916 15316
rect 27972 15260 29596 15316
rect 29652 15260 29662 15316
rect 31266 15260 31276 15316
rect 31332 15260 32956 15316
rect 33012 15260 33022 15316
rect 36082 15260 36092 15316
rect 36148 15260 37436 15316
rect 37492 15260 38220 15316
rect 38276 15260 38286 15316
rect 42354 15260 42364 15316
rect 42420 15260 43036 15316
rect 43092 15260 43102 15316
rect 45938 15260 45948 15316
rect 46004 15260 47068 15316
rect 47124 15260 47134 15316
rect 26852 15204 26908 15260
rect 7634 15148 7644 15204
rect 7700 15148 9548 15204
rect 9604 15148 9614 15204
rect 11890 15148 11900 15204
rect 11956 15148 11966 15204
rect 15708 15148 22428 15204
rect 22484 15148 22494 15204
rect 22754 15148 22764 15204
rect 22820 15148 24892 15204
rect 24948 15148 24958 15204
rect 25666 15148 25676 15204
rect 25732 15148 26460 15204
rect 26516 15148 26526 15204
rect 26852 15148 28364 15204
rect 28420 15148 28430 15204
rect 33394 15148 33404 15204
rect 33460 15148 33964 15204
rect 34020 15148 34030 15204
rect 51314 15148 51324 15204
rect 51380 15148 51884 15204
rect 51940 15148 51950 15204
rect 11900 15092 11956 15148
rect 11778 15036 11788 15092
rect 11844 15036 11956 15092
rect 15222 15036 15260 15092
rect 15316 15036 15326 15092
rect 20150 15036 20188 15092
rect 20244 15036 20254 15092
rect 20738 15036 20748 15092
rect 20804 15036 21084 15092
rect 21140 15036 21150 15092
rect 23538 15036 23548 15092
rect 23604 15036 25900 15092
rect 25956 15036 25966 15092
rect 30482 15036 30492 15092
rect 30548 15036 39228 15092
rect 39284 15036 39788 15092
rect 39844 15036 39854 15092
rect 40226 15036 40236 15092
rect 40292 15036 45612 15092
rect 45668 15036 45678 15092
rect 6626 14924 6636 14980
rect 6692 14924 8428 14980
rect 8484 14924 12908 14980
rect 12964 14924 12974 14980
rect 15474 14924 15484 14980
rect 15540 14924 22652 14980
rect 22708 14924 23660 14980
rect 23716 14924 23726 14980
rect 28102 14924 28140 14980
rect 28196 14924 28206 14980
rect 33394 14924 33404 14980
rect 33460 14924 33740 14980
rect 33796 14924 33806 14980
rect 38546 14924 38556 14980
rect 38612 14924 41132 14980
rect 41188 14924 41198 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 5842 14812 5852 14868
rect 5908 14812 13692 14868
rect 13748 14812 13758 14868
rect 19618 14812 19628 14868
rect 19684 14812 20188 14868
rect 20244 14812 20254 14868
rect 20738 14812 20748 14868
rect 20804 14812 21756 14868
rect 21812 14812 21822 14868
rect 22540 14812 25116 14868
rect 25172 14812 25182 14868
rect 31490 14812 31500 14868
rect 31556 14812 31836 14868
rect 31892 14812 31902 14868
rect 42130 14812 42140 14868
rect 42196 14812 43484 14868
rect 43540 14812 43550 14868
rect 45826 14812 45836 14868
rect 45892 14812 46620 14868
rect 46676 14812 46686 14868
rect 22540 14756 22596 14812
rect 10546 14700 10556 14756
rect 10612 14700 22596 14756
rect 22754 14700 22764 14756
rect 22820 14700 24108 14756
rect 24164 14700 25676 14756
rect 25732 14700 25742 14756
rect 33506 14700 33516 14756
rect 33572 14700 41132 14756
rect 41188 14700 42364 14756
rect 42420 14700 42430 14756
rect 5170 14588 5180 14644
rect 5236 14588 5852 14644
rect 5908 14588 5918 14644
rect 7186 14588 7196 14644
rect 7252 14588 7868 14644
rect 7924 14588 7934 14644
rect 8306 14588 8316 14644
rect 8372 14588 12684 14644
rect 12740 14588 13468 14644
rect 13524 14588 13534 14644
rect 14578 14588 14588 14644
rect 14644 14588 17500 14644
rect 17556 14588 17566 14644
rect 20626 14588 20636 14644
rect 20692 14588 26908 14644
rect 26964 14588 26974 14644
rect 32386 14588 32396 14644
rect 32452 14588 33628 14644
rect 33684 14588 33694 14644
rect 35522 14588 35532 14644
rect 35588 14588 36316 14644
rect 36372 14588 36382 14644
rect 38546 14588 38556 14644
rect 38612 14588 43148 14644
rect 43204 14588 43214 14644
rect 43810 14588 43820 14644
rect 43876 14588 46172 14644
rect 46228 14588 46396 14644
rect 46452 14588 46462 14644
rect 6178 14476 6188 14532
rect 6244 14476 12572 14532
rect 12628 14476 15260 14532
rect 15316 14476 15326 14532
rect 21186 14476 21196 14532
rect 21252 14476 21532 14532
rect 21588 14476 21598 14532
rect 23660 14476 32172 14532
rect 32228 14476 32238 14532
rect 35074 14476 35084 14532
rect 35140 14476 39004 14532
rect 39060 14476 39452 14532
rect 39508 14476 39518 14532
rect 53330 14476 53340 14532
rect 53396 14476 55580 14532
rect 55636 14476 55646 14532
rect 23660 14420 23716 14476
rect 5394 14364 5404 14420
rect 5460 14364 6524 14420
rect 6580 14364 8652 14420
rect 8708 14364 8718 14420
rect 10882 14364 10892 14420
rect 10948 14364 12124 14420
rect 12180 14364 12684 14420
rect 12740 14364 12750 14420
rect 15922 14364 15932 14420
rect 15988 14364 21084 14420
rect 21140 14364 21150 14420
rect 22306 14364 22316 14420
rect 22372 14364 23100 14420
rect 23156 14364 23166 14420
rect 23650 14364 23660 14420
rect 23716 14364 23726 14420
rect 26226 14364 26236 14420
rect 26292 14364 27132 14420
rect 27188 14364 27198 14420
rect 27794 14364 27804 14420
rect 27860 14364 29372 14420
rect 29428 14364 29438 14420
rect 31938 14364 31948 14420
rect 32004 14364 33628 14420
rect 33684 14364 34972 14420
rect 35028 14364 35038 14420
rect 38658 14364 38668 14420
rect 38724 14364 39116 14420
rect 39172 14364 39182 14420
rect 42802 14364 42812 14420
rect 42868 14364 45052 14420
rect 45108 14364 45118 14420
rect 7410 14252 7420 14308
rect 7476 14252 9324 14308
rect 9380 14252 9390 14308
rect 19282 14252 19292 14308
rect 19348 14252 19740 14308
rect 19796 14252 19806 14308
rect 20188 14252 25004 14308
rect 25060 14252 25070 14308
rect 28130 14252 28140 14308
rect 28196 14252 30492 14308
rect 30548 14252 30558 14308
rect 41794 14252 41804 14308
rect 41860 14252 43148 14308
rect 43204 14252 43214 14308
rect 44930 14252 44940 14308
rect 44996 14252 45724 14308
rect 45780 14252 45790 14308
rect 46162 14252 46172 14308
rect 46228 14252 47068 14308
rect 47124 14252 47134 14308
rect 14466 14140 14476 14196
rect 14532 14140 14924 14196
rect 14980 14140 14990 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 13682 14028 13692 14084
rect 13748 14028 19516 14084
rect 19572 14028 19582 14084
rect 20188 13972 20244 14252
rect 21298 14140 21308 14196
rect 21364 14140 24220 14196
rect 24276 14140 26572 14196
rect 26628 14140 26638 14196
rect 33282 14140 33292 14196
rect 33348 14140 35308 14196
rect 35364 14140 35374 14196
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 22194 14028 22204 14084
rect 22260 14028 23996 14084
rect 24052 14028 24062 14084
rect 30482 14028 30492 14084
rect 30548 14028 31276 14084
rect 31332 14028 31342 14084
rect 35084 14028 41468 14084
rect 41524 14028 42252 14084
rect 42308 14028 42318 14084
rect 7718 13916 7756 13972
rect 7812 13916 7822 13972
rect 8306 13916 8316 13972
rect 8372 13916 8876 13972
rect 8932 13916 8942 13972
rect 9090 13916 9100 13972
rect 9156 13916 11228 13972
rect 11284 13916 11294 13972
rect 11778 13916 11788 13972
rect 11844 13916 20244 13972
rect 20626 13916 20636 13972
rect 20692 13916 21532 13972
rect 21588 13916 21598 13972
rect 23286 13916 23324 13972
rect 23380 13916 23390 13972
rect 23538 13916 23548 13972
rect 23604 13916 23642 13972
rect 35084 13860 35140 14028
rect 39340 13916 43708 13972
rect 45154 13916 45164 13972
rect 45220 13916 46508 13972
rect 46564 13916 47404 13972
rect 47460 13916 47470 13972
rect 39340 13860 39396 13916
rect 43652 13860 43708 13916
rect 9996 13804 15148 13860
rect 16818 13804 16828 13860
rect 16884 13804 19180 13860
rect 19236 13804 19246 13860
rect 19730 13804 19740 13860
rect 19796 13804 22428 13860
rect 22484 13804 22494 13860
rect 23650 13804 23660 13860
rect 23716 13804 23772 13860
rect 23828 13804 23838 13860
rect 24770 13804 24780 13860
rect 24836 13804 29484 13860
rect 29540 13804 30492 13860
rect 30548 13804 30558 13860
rect 31042 13804 31052 13860
rect 31108 13804 33628 13860
rect 33684 13804 33694 13860
rect 35074 13804 35084 13860
rect 35140 13804 35150 13860
rect 37762 13804 37772 13860
rect 37828 13804 38892 13860
rect 38948 13804 38958 13860
rect 39330 13804 39340 13860
rect 39396 13804 39406 13860
rect 43474 13804 43484 13860
rect 43540 13804 43550 13860
rect 43652 13804 44828 13860
rect 44884 13804 44894 13860
rect 45490 13804 45500 13860
rect 45556 13804 46732 13860
rect 46788 13804 46798 13860
rect 9996 13748 10052 13804
rect 15092 13748 15148 13804
rect 43484 13748 43540 13804
rect 6626 13692 6636 13748
rect 6692 13692 10052 13748
rect 10210 13692 10220 13748
rect 10276 13692 11340 13748
rect 11396 13692 11406 13748
rect 11890 13692 11900 13748
rect 11956 13692 14924 13748
rect 14980 13692 14990 13748
rect 15092 13692 16268 13748
rect 16324 13692 18396 13748
rect 18452 13692 18462 13748
rect 18946 13692 18956 13748
rect 19012 13692 20636 13748
rect 20692 13692 20702 13748
rect 20850 13692 20860 13748
rect 20916 13692 20972 13748
rect 21028 13692 21038 13748
rect 22978 13692 22988 13748
rect 23044 13692 27804 13748
rect 27860 13692 27870 13748
rect 29362 13692 29372 13748
rect 29428 13692 30604 13748
rect 30660 13692 30670 13748
rect 32274 13692 32284 13748
rect 32340 13692 33852 13748
rect 33908 13692 35196 13748
rect 35252 13692 35262 13748
rect 37986 13692 37996 13748
rect 38052 13692 38668 13748
rect 38724 13692 38734 13748
rect 43484 13692 45836 13748
rect 45892 13692 45902 13748
rect 46386 13692 46396 13748
rect 46452 13692 47292 13748
rect 47348 13692 47358 13748
rect 49522 13692 49532 13748
rect 49588 13692 52220 13748
rect 52276 13692 52286 13748
rect 8194 13580 8204 13636
rect 8260 13580 10332 13636
rect 10388 13580 11004 13636
rect 11060 13580 11070 13636
rect 15362 13580 15372 13636
rect 15428 13580 16940 13636
rect 16996 13580 17006 13636
rect 18386 13580 18396 13636
rect 18452 13580 21868 13636
rect 21924 13580 21934 13636
rect 26338 13580 26348 13636
rect 26404 13580 28588 13636
rect 28644 13580 28654 13636
rect 29138 13580 29148 13636
rect 29204 13580 29932 13636
rect 29988 13580 29998 13636
rect 32498 13580 32508 13636
rect 32564 13580 34636 13636
rect 34692 13580 34702 13636
rect 43474 13580 43484 13636
rect 43540 13580 45388 13636
rect 45444 13580 46172 13636
rect 46228 13580 46238 13636
rect 59200 13524 60000 13552
rect 10210 13468 10220 13524
rect 10276 13468 10892 13524
rect 10948 13468 10958 13524
rect 16370 13468 16380 13524
rect 16436 13468 18060 13524
rect 18116 13468 18126 13524
rect 18498 13468 18508 13524
rect 18564 13468 18956 13524
rect 19012 13468 19022 13524
rect 20066 13468 20076 13524
rect 20132 13468 21420 13524
rect 21476 13468 21486 13524
rect 22754 13468 22764 13524
rect 22820 13468 23548 13524
rect 23604 13468 23614 13524
rect 25442 13468 25452 13524
rect 25508 13468 26684 13524
rect 26740 13468 26750 13524
rect 29586 13468 29596 13524
rect 29652 13468 29662 13524
rect 45602 13468 45612 13524
rect 45668 13468 47292 13524
rect 47348 13468 47358 13524
rect 58146 13468 58156 13524
rect 58212 13468 60000 13524
rect 29596 13412 29652 13468
rect 59200 13440 60000 13468
rect 7830 13356 7868 13412
rect 7924 13356 7934 13412
rect 14028 13356 27692 13412
rect 27748 13356 27758 13412
rect 28914 13356 28924 13412
rect 28980 13356 29652 13412
rect 41906 13356 41916 13412
rect 41972 13356 43036 13412
rect 43092 13356 43102 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 6178 13020 6188 13076
rect 6244 13020 10108 13076
rect 10164 13020 10174 13076
rect 12898 13020 12908 13076
rect 12964 13020 13244 13076
rect 13300 13020 13310 13076
rect 14028 12964 14084 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 22726 13244 22764 13300
rect 22820 13244 22830 13300
rect 23090 13244 23100 13300
rect 23156 13244 23884 13300
rect 23940 13244 23950 13300
rect 24108 13244 26908 13300
rect 26964 13244 26974 13300
rect 24108 13188 24164 13244
rect 15026 13132 15036 13188
rect 15092 13132 15148 13188
rect 15204 13132 15596 13188
rect 15652 13132 15662 13188
rect 18386 13132 18396 13188
rect 18452 13132 24164 13188
rect 25078 13132 25116 13188
rect 25172 13132 25182 13188
rect 27234 13132 27244 13188
rect 27300 13132 28476 13188
rect 28532 13132 28542 13188
rect 20178 13020 20188 13076
rect 20244 13020 20804 13076
rect 24182 13020 24220 13076
rect 24276 13020 24286 13076
rect 25666 13020 25676 13076
rect 25732 13020 27916 13076
rect 27972 13020 27982 13076
rect 46834 13020 46844 13076
rect 46900 13020 48972 13076
rect 49028 13020 50092 13076
rect 50148 13020 50158 13076
rect 20748 12964 20804 13020
rect 6962 12908 6972 12964
rect 7028 12908 14028 12964
rect 14084 12908 14094 12964
rect 20738 12908 20748 12964
rect 20804 12908 20814 12964
rect 22390 12908 22428 12964
rect 22484 12908 22494 12964
rect 27682 12908 27692 12964
rect 27748 12908 28140 12964
rect 28196 12908 28206 12964
rect 42018 12908 42028 12964
rect 42084 12908 42588 12964
rect 42644 12908 42654 12964
rect 49186 12908 49196 12964
rect 49252 12908 50204 12964
rect 50260 12908 50270 12964
rect 6738 12796 6748 12852
rect 6804 12796 7308 12852
rect 7364 12796 8652 12852
rect 8708 12796 12348 12852
rect 12404 12796 14588 12852
rect 14644 12796 14654 12852
rect 17574 12796 17612 12852
rect 17668 12796 17678 12852
rect 13682 12684 13692 12740
rect 13748 12684 15148 12740
rect 16594 12684 16604 12740
rect 16660 12684 27692 12740
rect 27748 12684 27758 12740
rect 31042 12684 31052 12740
rect 31108 12684 31388 12740
rect 31444 12684 31454 12740
rect 15092 12628 15148 12684
rect 15092 12572 15932 12628
rect 15988 12572 15998 12628
rect 21970 12572 21980 12628
rect 22036 12572 22876 12628
rect 22932 12572 22942 12628
rect 28130 12572 28140 12628
rect 28196 12572 31500 12628
rect 31556 12572 31566 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 12002 12460 12012 12516
rect 12068 12460 15372 12516
rect 15428 12460 15438 12516
rect 16370 12460 16380 12516
rect 16436 12460 18116 12516
rect 24434 12460 24444 12516
rect 24500 12460 25564 12516
rect 25620 12460 25630 12516
rect 27346 12460 27356 12516
rect 27412 12460 28140 12516
rect 28196 12460 28206 12516
rect 30716 12460 31052 12516
rect 31108 12460 31118 12516
rect 18060 12404 18116 12460
rect 30716 12404 30772 12460
rect 7298 12348 7308 12404
rect 7364 12348 8204 12404
rect 8260 12348 8270 12404
rect 9650 12348 9660 12404
rect 9716 12348 11228 12404
rect 11284 12348 15260 12404
rect 15316 12348 17052 12404
rect 17108 12348 17118 12404
rect 17490 12348 17500 12404
rect 17556 12348 17566 12404
rect 17798 12348 17836 12404
rect 17892 12348 17902 12404
rect 18060 12348 30772 12404
rect 30930 12348 30940 12404
rect 30996 12348 31388 12404
rect 31444 12348 35196 12404
rect 35252 12348 35756 12404
rect 35812 12348 36428 12404
rect 36484 12348 36876 12404
rect 36932 12348 36942 12404
rect 10210 12236 10220 12292
rect 10276 12236 11900 12292
rect 11956 12236 11966 12292
rect 17500 12180 17556 12348
rect 20402 12236 20412 12292
rect 20468 12236 26124 12292
rect 26180 12236 27580 12292
rect 27636 12236 27646 12292
rect 27804 12236 30044 12292
rect 30100 12236 30110 12292
rect 30258 12236 30268 12292
rect 30324 12236 31108 12292
rect 47506 12236 47516 12292
rect 47572 12236 49196 12292
rect 49252 12236 49262 12292
rect 27804 12180 27860 12236
rect 31052 12180 31108 12236
rect 59200 12180 60000 12208
rect 8754 12124 8764 12180
rect 8820 12124 11340 12180
rect 11396 12124 11406 12180
rect 11666 12124 11676 12180
rect 11732 12124 16268 12180
rect 16324 12124 17556 12180
rect 18946 12124 18956 12180
rect 19012 12124 21308 12180
rect 21364 12124 21374 12180
rect 21746 12124 21756 12180
rect 21812 12124 22428 12180
rect 22484 12124 22494 12180
rect 22642 12124 22652 12180
rect 22708 12124 23212 12180
rect 23268 12124 27356 12180
rect 27412 12124 27422 12180
rect 27570 12124 27580 12180
rect 27636 12124 27646 12180
rect 27794 12124 27804 12180
rect 27860 12124 27870 12180
rect 29922 12124 29932 12180
rect 29988 12124 30492 12180
rect 30548 12124 30558 12180
rect 31042 12124 31052 12180
rect 31108 12124 34748 12180
rect 34804 12124 35980 12180
rect 36036 12124 36046 12180
rect 42914 12124 42924 12180
rect 42980 12124 43372 12180
rect 43428 12124 44492 12180
rect 44548 12124 44558 12180
rect 58146 12124 58156 12180
rect 58212 12124 60000 12180
rect 27580 12068 27636 12124
rect 59200 12096 60000 12124
rect 10770 12012 10780 12068
rect 10836 12012 11788 12068
rect 11844 12012 14028 12068
rect 14084 12012 14094 12068
rect 15092 12012 27356 12068
rect 27412 12012 27422 12068
rect 27580 12012 29260 12068
rect 29316 12012 29708 12068
rect 29764 12012 29774 12068
rect 41682 12012 41692 12068
rect 41748 12012 42588 12068
rect 42644 12012 42654 12068
rect 44034 12012 44044 12068
rect 44100 12012 46620 12068
rect 46676 12012 46686 12068
rect 7858 11900 7868 11956
rect 7924 11900 13412 11956
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 13356 11732 13412 11900
rect 15092 11844 15148 12012
rect 16706 11900 16716 11956
rect 16772 11900 18956 11956
rect 19012 11900 19022 11956
rect 20178 11900 20188 11956
rect 20244 11900 21980 11956
rect 22036 11900 22652 11956
rect 22708 11900 22718 11956
rect 22866 11900 22876 11956
rect 22932 11900 22970 11956
rect 24210 11900 24220 11956
rect 24276 11900 24556 11956
rect 24612 11900 24622 11956
rect 26898 11900 26908 11956
rect 26964 11900 28700 11956
rect 28756 11900 28766 11956
rect 31154 11900 31164 11956
rect 31220 11900 35868 11956
rect 35924 11900 35934 11956
rect 13570 11788 13580 11844
rect 13636 11788 15148 11844
rect 15474 11788 15484 11844
rect 15540 11788 16940 11844
rect 16996 11788 17006 11844
rect 17154 11788 17164 11844
rect 17220 11788 17500 11844
rect 17556 11788 17566 11844
rect 19170 11788 19180 11844
rect 19236 11788 20860 11844
rect 20916 11788 20926 11844
rect 21830 11788 21868 11844
rect 21924 11788 21934 11844
rect 23762 11788 23772 11844
rect 23828 11788 25116 11844
rect 25172 11788 25788 11844
rect 25844 11788 26572 11844
rect 26628 11788 26638 11844
rect 27346 11788 27356 11844
rect 27412 11788 28812 11844
rect 28868 11788 28878 11844
rect 36950 11788 36988 11844
rect 37044 11788 37054 11844
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 7522 11676 7532 11732
rect 7588 11676 8316 11732
rect 8372 11676 8382 11732
rect 10434 11676 10444 11732
rect 10500 11676 12796 11732
rect 12852 11676 12862 11732
rect 13356 11676 16156 11732
rect 16212 11676 16222 11732
rect 16706 11676 16716 11732
rect 16772 11676 20748 11732
rect 20804 11676 20814 11732
rect 24322 11676 24332 11732
rect 24388 11676 24892 11732
rect 24948 11676 24958 11732
rect 27234 11676 27244 11732
rect 27300 11676 28476 11732
rect 28532 11676 30156 11732
rect 30212 11676 30222 11732
rect 36082 11676 36092 11732
rect 36148 11676 38780 11732
rect 38836 11676 38846 11732
rect 10444 11620 10500 11676
rect 6626 11564 6636 11620
rect 6692 11564 7756 11620
rect 7812 11564 10500 11620
rect 11218 11564 11228 11620
rect 11284 11564 11900 11620
rect 11956 11564 13580 11620
rect 13636 11564 13646 11620
rect 15698 11564 15708 11620
rect 15764 11564 22540 11620
rect 22596 11564 22606 11620
rect 22978 11564 22988 11620
rect 23044 11564 23436 11620
rect 23492 11564 23502 11620
rect 24322 11564 24332 11620
rect 24388 11564 25004 11620
rect 25060 11564 25070 11620
rect 25442 11564 25452 11620
rect 25508 11564 25900 11620
rect 25956 11564 25966 11620
rect 32946 11564 32956 11620
rect 33012 11564 33740 11620
rect 33796 11564 33806 11620
rect 34178 11564 34188 11620
rect 34244 11564 36652 11620
rect 36708 11564 37324 11620
rect 37380 11564 37390 11620
rect 11228 11508 11284 11564
rect 59200 11508 60000 11536
rect 7074 11452 7084 11508
rect 7140 11452 11284 11508
rect 16930 11452 16940 11508
rect 16996 11452 18228 11508
rect 18358 11452 18396 11508
rect 18452 11452 18462 11508
rect 18610 11452 18620 11508
rect 18676 11452 25676 11508
rect 25732 11452 27244 11508
rect 27300 11452 27310 11508
rect 28690 11452 28700 11508
rect 28756 11452 29596 11508
rect 29652 11452 29662 11508
rect 31378 11452 31388 11508
rect 31444 11452 34300 11508
rect 34356 11452 34748 11508
rect 34804 11452 34814 11508
rect 35186 11452 35196 11508
rect 35252 11452 36092 11508
rect 36148 11452 36158 11508
rect 40338 11452 40348 11508
rect 40404 11452 41132 11508
rect 41188 11452 41198 11508
rect 57922 11452 57932 11508
rect 57988 11452 60000 11508
rect 18172 11396 18228 11452
rect 59200 11424 60000 11452
rect 8082 11340 8092 11396
rect 8148 11340 9212 11396
rect 9268 11340 9278 11396
rect 9762 11340 9772 11396
rect 9828 11340 10220 11396
rect 10276 11340 11900 11396
rect 11956 11340 11966 11396
rect 15026 11340 15036 11396
rect 15092 11340 17388 11396
rect 17444 11340 17454 11396
rect 18172 11340 22932 11396
rect 23090 11340 23100 11396
rect 23156 11340 23772 11396
rect 23828 11340 23838 11396
rect 24070 11340 24108 11396
rect 24164 11340 24174 11396
rect 24546 11340 24556 11396
rect 24612 11340 26572 11396
rect 26628 11340 26638 11396
rect 28802 11340 28812 11396
rect 28868 11340 31052 11396
rect 31108 11340 31118 11396
rect 33506 11340 33516 11396
rect 33572 11340 34076 11396
rect 34132 11340 34142 11396
rect 34626 11340 34636 11396
rect 34692 11340 35308 11396
rect 35364 11340 35374 11396
rect 38612 11340 39452 11396
rect 39508 11340 40460 11396
rect 40516 11340 40526 11396
rect 41794 11340 41804 11396
rect 41860 11340 42028 11396
rect 42084 11340 43372 11396
rect 43428 11340 43708 11396
rect 43764 11340 43774 11396
rect 46946 11340 46956 11396
rect 47012 11340 47516 11396
rect 47572 11340 47582 11396
rect 51650 11340 51660 11396
rect 51716 11340 55580 11396
rect 55636 11340 55646 11396
rect 22876 11284 22932 11340
rect 38612 11284 38668 11340
rect 12338 11228 12348 11284
rect 12404 11228 15820 11284
rect 15876 11228 16716 11284
rect 16772 11228 16782 11284
rect 17154 11228 17164 11284
rect 17220 11228 18172 11284
rect 18228 11228 19516 11284
rect 19572 11228 21364 11284
rect 22876 11228 25452 11284
rect 25508 11228 25518 11284
rect 29250 11228 29260 11284
rect 29316 11228 29932 11284
rect 29988 11228 30940 11284
rect 30996 11228 31006 11284
rect 34514 11228 34524 11284
rect 34580 11228 38668 11284
rect 42242 11228 42252 11284
rect 42308 11228 43932 11284
rect 43988 11228 43998 11284
rect 10098 11116 10108 11172
rect 10164 11116 12908 11172
rect 12964 11116 12974 11172
rect 15092 11116 19404 11172
rect 19460 11116 19852 11172
rect 19908 11116 19918 11172
rect 20178 11116 20188 11172
rect 20244 11116 21084 11172
rect 21140 11116 21150 11172
rect 15092 11060 15148 11116
rect 8754 11004 8764 11060
rect 8820 11004 14028 11060
rect 14084 11004 15148 11060
rect 16492 11004 16940 11060
rect 16996 11004 17006 11060
rect 16492 10948 16548 11004
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 21308 10948 21364 11228
rect 23874 11116 23884 11172
rect 23940 11116 24332 11172
rect 24388 11116 24398 11172
rect 24546 11116 24556 11172
rect 24612 11116 24650 11172
rect 25778 11116 25788 11172
rect 25844 11116 27412 11172
rect 27570 11116 27580 11172
rect 27636 11116 38668 11172
rect 41682 11116 41692 11172
rect 41748 11116 42924 11172
rect 42980 11116 42990 11172
rect 47842 11116 47852 11172
rect 47908 11116 48972 11172
rect 49028 11116 49038 11172
rect 27356 11060 27412 11116
rect 21746 11004 21756 11060
rect 21812 11004 27020 11060
rect 27076 11004 27086 11060
rect 27356 11004 33796 11060
rect 33740 10948 33796 11004
rect 38612 10948 38668 11116
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 8204 10892 10556 10948
rect 10612 10892 10622 10948
rect 12786 10892 12796 10948
rect 12852 10892 16548 10948
rect 16604 10892 18508 10948
rect 18564 10892 18574 10948
rect 21308 10892 24164 10948
rect 33730 10892 33740 10948
rect 33796 10892 33806 10948
rect 38612 10892 42140 10948
rect 42196 10892 42206 10948
rect 8204 10836 8260 10892
rect 16604 10836 16660 10892
rect 24108 10836 24164 10892
rect 59200 10836 60000 10864
rect 7410 10780 7420 10836
rect 7476 10780 8204 10836
rect 8260 10780 8270 10836
rect 10434 10780 10444 10836
rect 10500 10780 12572 10836
rect 12628 10780 12638 10836
rect 12898 10780 12908 10836
rect 12964 10780 16660 10836
rect 16818 10780 16828 10836
rect 16884 10780 18172 10836
rect 18228 10780 18238 10836
rect 19058 10780 19068 10836
rect 19124 10780 19740 10836
rect 19796 10780 19806 10836
rect 22950 10780 22988 10836
rect 23044 10780 23054 10836
rect 24098 10780 24108 10836
rect 24164 10780 24174 10836
rect 24322 10780 24332 10836
rect 24388 10780 25004 10836
rect 25060 10780 25340 10836
rect 25396 10780 25406 10836
rect 30146 10780 30156 10836
rect 30212 10780 41468 10836
rect 41524 10780 41534 10836
rect 58146 10780 58156 10836
rect 58212 10780 60000 10836
rect 16604 10724 16660 10780
rect 59200 10752 60000 10780
rect 9090 10668 9100 10724
rect 9156 10668 15596 10724
rect 15652 10668 15662 10724
rect 16604 10668 16940 10724
rect 16996 10668 17006 10724
rect 18022 10668 18060 10724
rect 18116 10668 18126 10724
rect 19394 10668 19404 10724
rect 19460 10668 19628 10724
rect 19684 10668 19694 10724
rect 22530 10668 22540 10724
rect 22596 10668 22606 10724
rect 23734 10668 23772 10724
rect 23828 10668 23838 10724
rect 25330 10668 25340 10724
rect 25396 10668 25406 10724
rect 25750 10668 25788 10724
rect 25844 10668 25854 10724
rect 30594 10668 30604 10724
rect 30660 10668 31836 10724
rect 31892 10668 31902 10724
rect 33618 10668 33628 10724
rect 33684 10668 34972 10724
rect 35028 10668 39788 10724
rect 39844 10668 39854 10724
rect 11442 10556 11452 10612
rect 11508 10556 12348 10612
rect 12404 10556 13580 10612
rect 13636 10556 13646 10612
rect 16146 10556 16156 10612
rect 16212 10556 18956 10612
rect 19012 10556 19022 10612
rect 19506 10556 19516 10612
rect 19572 10556 20524 10612
rect 20580 10556 20590 10612
rect 10546 10444 10556 10500
rect 10612 10444 13468 10500
rect 13524 10444 18396 10500
rect 18452 10444 18462 10500
rect 19516 10388 19572 10556
rect 22540 10500 22596 10668
rect 25340 10612 25396 10668
rect 25340 10556 25676 10612
rect 25732 10556 25742 10612
rect 26002 10556 26012 10612
rect 26068 10556 26348 10612
rect 26404 10556 26414 10612
rect 33516 10556 35980 10612
rect 36036 10556 36046 10612
rect 37202 10556 37212 10612
rect 37268 10556 42364 10612
rect 42420 10556 42430 10612
rect 43026 10556 43036 10612
rect 43092 10556 46732 10612
rect 46788 10556 47180 10612
rect 47236 10556 47246 10612
rect 47618 10556 47628 10612
rect 47684 10556 48860 10612
rect 48916 10556 48926 10612
rect 22540 10444 26908 10500
rect 26964 10444 26974 10500
rect 29110 10444 29148 10500
rect 29204 10444 29214 10500
rect 30034 10444 30044 10500
rect 30100 10444 31276 10500
rect 31332 10444 31342 10500
rect 15362 10332 15372 10388
rect 15428 10332 15708 10388
rect 15764 10332 15774 10388
rect 18050 10332 18060 10388
rect 18116 10332 19572 10388
rect 21074 10332 21084 10388
rect 21140 10332 22764 10388
rect 22820 10332 22830 10388
rect 23090 10332 23100 10388
rect 23156 10332 29932 10388
rect 29988 10332 29998 10388
rect 18386 10220 18396 10276
rect 18452 10220 32956 10276
rect 33012 10220 33022 10276
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 33516 10164 33572 10556
rect 35980 10500 36036 10556
rect 35980 10444 37548 10500
rect 37604 10444 37614 10500
rect 38612 10444 39676 10500
rect 39732 10444 39742 10500
rect 38612 10388 38668 10444
rect 34066 10332 34076 10388
rect 34132 10332 35420 10388
rect 35476 10332 37884 10388
rect 37940 10332 38668 10388
rect 38546 10220 38556 10276
rect 38612 10220 39340 10276
rect 39396 10220 39406 10276
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 59200 10164 60000 10192
rect 19254 10108 19292 10164
rect 19348 10108 19358 10164
rect 20290 10108 20300 10164
rect 20356 10108 22092 10164
rect 22148 10108 23436 10164
rect 23492 10108 23502 10164
rect 24434 10108 24444 10164
rect 24500 10108 33572 10164
rect 57698 10108 57708 10164
rect 57764 10108 60000 10164
rect 59200 10080 60000 10108
rect 11638 9996 11676 10052
rect 11732 9996 11742 10052
rect 14914 9996 14924 10052
rect 14980 9996 20748 10052
rect 20804 9996 21644 10052
rect 21700 9996 21710 10052
rect 23314 9996 23324 10052
rect 23380 9996 24108 10052
rect 24164 9996 24174 10052
rect 24994 9996 25004 10052
rect 25060 9996 25452 10052
rect 25508 9996 27580 10052
rect 27636 9996 27646 10052
rect 30258 9996 30268 10052
rect 30324 9996 31724 10052
rect 31780 9996 31790 10052
rect 32610 9996 32620 10052
rect 32676 9996 36988 10052
rect 37044 9996 37054 10052
rect 40450 9996 40460 10052
rect 40516 9996 45388 10052
rect 45444 9996 45454 10052
rect 9426 9884 9436 9940
rect 9492 9884 12796 9940
rect 12852 9884 12862 9940
rect 14662 9884 14700 9940
rect 14756 9884 14766 9940
rect 16716 9884 19964 9940
rect 20020 9884 20030 9940
rect 21746 9884 21756 9940
rect 21812 9884 27468 9940
rect 27524 9884 27534 9940
rect 35858 9884 35868 9940
rect 35924 9884 37212 9940
rect 37268 9884 37278 9940
rect 46274 9884 46284 9940
rect 46340 9884 47068 9940
rect 47124 9884 47134 9940
rect 10322 9772 10332 9828
rect 10388 9772 12236 9828
rect 12292 9772 12302 9828
rect 13794 9772 13804 9828
rect 13860 9772 14252 9828
rect 14308 9772 15148 9828
rect 15092 9716 15148 9772
rect 16716 9716 16772 9884
rect 17042 9772 17052 9828
rect 17108 9772 18060 9828
rect 18116 9772 18126 9828
rect 18610 9772 18620 9828
rect 18676 9772 19292 9828
rect 19348 9772 19358 9828
rect 20626 9772 20636 9828
rect 20692 9772 24220 9828
rect 24276 9772 24286 9828
rect 27682 9772 27692 9828
rect 27748 9772 28364 9828
rect 28420 9772 29148 9828
rect 29204 9772 29214 9828
rect 32956 9772 38668 9828
rect 38724 9772 38734 9828
rect 40002 9772 40012 9828
rect 40068 9772 43820 9828
rect 43876 9772 43886 9828
rect 44146 9772 44156 9828
rect 44212 9772 45052 9828
rect 45108 9772 45118 9828
rect 45378 9772 45388 9828
rect 45444 9772 46508 9828
rect 46564 9772 46574 9828
rect 8978 9660 8988 9716
rect 9044 9660 13692 9716
rect 13748 9660 13758 9716
rect 14812 9660 16772 9716
rect 18386 9660 18396 9716
rect 18452 9660 19236 9716
rect 19618 9660 19628 9716
rect 19684 9660 20524 9716
rect 20580 9660 20590 9716
rect 21074 9660 21084 9716
rect 21140 9660 22540 9716
rect 22596 9660 22606 9716
rect 25330 9660 25340 9716
rect 25396 9660 26572 9716
rect 26628 9660 26638 9716
rect 14812 9380 14868 9660
rect 19180 9604 19236 9660
rect 15922 9548 15932 9604
rect 15988 9548 17276 9604
rect 17332 9548 17342 9604
rect 18162 9548 18172 9604
rect 18228 9548 18620 9604
rect 18676 9548 18686 9604
rect 19170 9548 19180 9604
rect 19236 9548 19246 9604
rect 19366 9548 19404 9604
rect 19460 9548 19470 9604
rect 19628 9548 19740 9604
rect 19796 9548 19806 9604
rect 19954 9548 19964 9604
rect 20020 9548 20748 9604
rect 20804 9548 21980 9604
rect 22036 9548 22046 9604
rect 22642 9548 22652 9604
rect 22708 9548 31612 9604
rect 31668 9548 31678 9604
rect 19628 9492 19684 9548
rect 16706 9436 16716 9492
rect 16772 9436 18396 9492
rect 18452 9436 18462 9492
rect 18834 9436 18844 9492
rect 18900 9436 19684 9492
rect 22418 9436 22428 9492
rect 22484 9436 22764 9492
rect 22820 9436 22830 9492
rect 23762 9436 23772 9492
rect 23828 9436 29596 9492
rect 29652 9436 29662 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 32956 9380 33012 9772
rect 38546 9660 38556 9716
rect 38612 9660 40684 9716
rect 40740 9660 40750 9716
rect 41346 9660 41356 9716
rect 41412 9660 42588 9716
rect 42644 9660 42654 9716
rect 49074 9548 49084 9604
rect 49140 9548 49980 9604
rect 50036 9548 51436 9604
rect 51492 9548 51502 9604
rect 59200 9492 60000 9520
rect 58146 9436 58156 9492
rect 58212 9436 60000 9492
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 59200 9408 60000 9436
rect 9986 9324 9996 9380
rect 10052 9324 11116 9380
rect 11172 9324 14476 9380
rect 14532 9324 14542 9380
rect 14802 9324 14812 9380
rect 14868 9324 14878 9380
rect 15698 9324 15708 9380
rect 15764 9324 18732 9380
rect 18788 9324 18798 9380
rect 24098 9324 24108 9380
rect 24164 9324 24332 9380
rect 24388 9324 24398 9380
rect 25778 9324 25788 9380
rect 25844 9324 26460 9380
rect 26516 9324 27076 9380
rect 27346 9324 27356 9380
rect 27412 9324 33012 9380
rect 27020 9268 27076 9324
rect 10882 9212 10892 9268
rect 10948 9212 13468 9268
rect 13524 9212 13534 9268
rect 14354 9212 14364 9268
rect 14420 9212 15484 9268
rect 15540 9212 15550 9268
rect 15810 9212 15820 9268
rect 15876 9212 16940 9268
rect 16996 9212 17006 9268
rect 18946 9212 18956 9268
rect 19012 9212 19180 9268
rect 19236 9212 25956 9268
rect 26086 9212 26124 9268
rect 26180 9212 26190 9268
rect 26562 9212 26572 9268
rect 26628 9212 26796 9268
rect 26852 9212 26862 9268
rect 27020 9212 27916 9268
rect 27972 9212 29372 9268
rect 29428 9212 29438 9268
rect 31490 9212 31500 9268
rect 31556 9212 32396 9268
rect 32452 9212 36092 9268
rect 36148 9212 36764 9268
rect 36820 9212 37100 9268
rect 37156 9212 37166 9268
rect 39778 9212 39788 9268
rect 39844 9212 40460 9268
rect 40516 9212 40526 9268
rect 13906 9100 13916 9156
rect 13972 9100 14924 9156
rect 14980 9100 14990 9156
rect 15922 9100 15932 9156
rect 15988 9100 23884 9156
rect 23940 9100 23950 9156
rect 24098 9100 24108 9156
rect 24164 9100 24556 9156
rect 24612 9100 24622 9156
rect 10434 8988 10444 9044
rect 10500 8988 16156 9044
rect 16212 8988 16828 9044
rect 16884 8988 16894 9044
rect 19058 8988 19068 9044
rect 19124 8988 24444 9044
rect 24500 8988 24510 9044
rect 24770 8988 24780 9044
rect 24836 8988 25676 9044
rect 25732 8988 25742 9044
rect 25900 8932 25956 9212
rect 26562 9100 26572 9156
rect 26628 9100 29260 9156
rect 29316 9100 29708 9156
rect 29764 9100 29774 9156
rect 47842 9100 47852 9156
rect 47908 9100 49084 9156
rect 49140 9100 49150 9156
rect 43810 8988 43820 9044
rect 43876 8988 44940 9044
rect 44996 8988 45006 9044
rect 49522 8988 49532 9044
rect 49588 8988 50204 9044
rect 50260 8988 50652 9044
rect 50708 8988 50718 9044
rect 11330 8876 11340 8932
rect 11396 8876 11406 8932
rect 11666 8876 11676 8932
rect 11732 8876 12236 8932
rect 12292 8876 12302 8932
rect 12674 8876 12684 8932
rect 12740 8876 19124 8932
rect 19394 8876 19404 8932
rect 19460 8876 20524 8932
rect 20580 8876 20590 8932
rect 21634 8876 21644 8932
rect 21700 8876 23324 8932
rect 23380 8876 23390 8932
rect 25900 8876 27804 8932
rect 27860 8876 27870 8932
rect 32498 8876 32508 8932
rect 32564 8876 43708 8932
rect 48178 8876 48188 8932
rect 48244 8876 49196 8932
rect 49252 8876 49262 8932
rect 11340 8820 11396 8876
rect 19068 8820 19124 8876
rect 43652 8820 43708 8876
rect 59200 8820 60000 8848
rect 11340 8764 15820 8820
rect 15876 8764 18172 8820
rect 18228 8764 18620 8820
rect 18676 8764 18686 8820
rect 19068 8764 20188 8820
rect 20244 8764 20254 8820
rect 23090 8764 23100 8820
rect 23156 8764 26684 8820
rect 26740 8764 26750 8820
rect 43652 8764 44268 8820
rect 44324 8764 44716 8820
rect 44772 8764 44782 8820
rect 59052 8764 60000 8820
rect 11330 8652 11340 8708
rect 11396 8652 12348 8708
rect 12404 8652 12414 8708
rect 15586 8652 15596 8708
rect 15652 8652 16996 8708
rect 17154 8652 17164 8708
rect 17220 8652 17612 8708
rect 17668 8652 17678 8708
rect 18386 8652 18396 8708
rect 18452 8652 25340 8708
rect 25396 8652 26012 8708
rect 26068 8652 26796 8708
rect 26852 8652 26862 8708
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 16940 8596 16996 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 13010 8540 13020 8596
rect 13076 8540 15708 8596
rect 15764 8540 16492 8596
rect 16548 8540 16558 8596
rect 16940 8540 18508 8596
rect 18564 8540 21084 8596
rect 21140 8540 22428 8596
rect 22484 8540 22494 8596
rect 25778 8540 25788 8596
rect 25844 8540 32004 8596
rect 13458 8428 13468 8484
rect 13524 8428 18732 8484
rect 18788 8428 19180 8484
rect 19236 8428 19246 8484
rect 19590 8428 19628 8484
rect 19684 8428 19694 8484
rect 20178 8428 20188 8484
rect 20244 8428 21980 8484
rect 22036 8428 22046 8484
rect 22306 8428 22316 8484
rect 22372 8428 23324 8484
rect 23380 8428 23390 8484
rect 24994 8428 25004 8484
rect 25060 8428 30268 8484
rect 30324 8428 30334 8484
rect 31948 8372 32004 8540
rect 59052 8484 59108 8764
rect 59200 8736 60000 8764
rect 59052 8428 59332 8484
rect 59276 8372 59332 8428
rect 14018 8316 14028 8372
rect 14084 8316 14924 8372
rect 14980 8316 14990 8372
rect 15922 8316 15932 8372
rect 15988 8316 16380 8372
rect 16436 8316 16716 8372
rect 16772 8316 16782 8372
rect 17500 8316 21420 8372
rect 21476 8316 21486 8372
rect 24882 8316 24892 8372
rect 24948 8316 25228 8372
rect 25284 8316 25294 8372
rect 31948 8316 35308 8372
rect 35364 8316 35374 8372
rect 42802 8316 42812 8372
rect 42868 8316 42878 8372
rect 43138 8316 43148 8372
rect 43204 8316 43708 8372
rect 43764 8316 43774 8372
rect 43922 8316 43932 8372
rect 43988 8316 45388 8372
rect 45444 8316 45454 8372
rect 57922 8316 57932 8372
rect 57988 8316 59332 8372
rect 9874 8204 9884 8260
rect 9940 8204 13804 8260
rect 13860 8204 13870 8260
rect 14354 8204 14364 8260
rect 14420 8204 15036 8260
rect 15092 8204 15372 8260
rect 15428 8204 15438 8260
rect 13804 8148 13860 8204
rect 15932 8148 15988 8316
rect 16258 8204 16268 8260
rect 16324 8204 16828 8260
rect 16884 8204 16894 8260
rect 17500 8148 17556 8316
rect 42812 8260 42868 8316
rect 18162 8204 18172 8260
rect 18228 8204 26908 8260
rect 31714 8204 31724 8260
rect 31780 8204 32060 8260
rect 32116 8204 32126 8260
rect 41458 8204 41468 8260
rect 41524 8204 42476 8260
rect 42532 8204 42868 8260
rect 43026 8204 43036 8260
rect 43092 8204 45164 8260
rect 45220 8204 45230 8260
rect 45490 8204 45500 8260
rect 45556 8204 45566 8260
rect 51986 8204 51996 8260
rect 52052 8204 55580 8260
rect 55636 8204 55646 8260
rect 26852 8148 26908 8204
rect 45500 8148 45556 8204
rect 59200 8148 60000 8176
rect 12002 8092 12012 8148
rect 12068 8092 13356 8148
rect 13412 8092 13422 8148
rect 13804 8092 15988 8148
rect 16146 8092 16156 8148
rect 16212 8092 17388 8148
rect 17444 8092 17556 8148
rect 18386 8092 18396 8148
rect 18452 8092 19964 8148
rect 20020 8092 20030 8148
rect 21522 8092 21532 8148
rect 21588 8092 23772 8148
rect 23828 8092 23838 8148
rect 24994 8092 25004 8148
rect 25060 8092 25788 8148
rect 25844 8092 25854 8148
rect 26852 8092 27580 8148
rect 27636 8092 27646 8148
rect 28354 8092 28364 8148
rect 28420 8092 30044 8148
rect 30100 8092 30110 8148
rect 30370 8092 30380 8148
rect 30436 8092 33068 8148
rect 33124 8092 33134 8148
rect 36082 8092 36092 8148
rect 36148 8092 38668 8148
rect 43698 8092 43708 8148
rect 43764 8092 45556 8148
rect 58146 8092 58156 8148
rect 58212 8092 60000 8148
rect 15362 7980 15372 8036
rect 15428 7980 21868 8036
rect 21924 7980 21934 8036
rect 26310 7980 26348 8036
rect 26404 7980 26414 8036
rect 27234 7980 27244 8036
rect 27300 7980 28476 8036
rect 28532 7980 28542 8036
rect 29586 7980 29596 8036
rect 29652 7980 30156 8036
rect 30212 7980 30222 8036
rect 32050 7980 32060 8036
rect 32116 7980 32732 8036
rect 32788 7980 33180 8036
rect 33236 7980 35532 8036
rect 35588 7980 35598 8036
rect 38612 7924 38668 8092
rect 59200 8064 60000 8092
rect 39106 7980 39116 8036
rect 39172 7980 43372 8036
rect 43428 7980 43438 8036
rect 15250 7868 15260 7924
rect 15316 7868 18172 7924
rect 18228 7868 18238 7924
rect 22866 7868 22876 7924
rect 22932 7868 23660 7924
rect 23716 7868 24556 7924
rect 24612 7868 24622 7924
rect 38612 7868 45500 7924
rect 45556 7868 46172 7924
rect 46228 7868 46238 7924
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 20934 7756 20972 7812
rect 21028 7756 21038 7812
rect 32508 7756 42700 7812
rect 42756 7756 42766 7812
rect 15474 7644 15484 7700
rect 15540 7644 15932 7700
rect 15988 7644 17948 7700
rect 18004 7644 20076 7700
rect 20132 7644 20142 7700
rect 20374 7644 20412 7700
rect 20468 7644 20478 7700
rect 20626 7644 20636 7700
rect 20692 7644 21868 7700
rect 21924 7644 21934 7700
rect 23874 7644 23884 7700
rect 23940 7644 25788 7700
rect 25844 7644 25854 7700
rect 28242 7644 28252 7700
rect 28308 7644 29036 7700
rect 29092 7644 29102 7700
rect 20636 7588 20692 7644
rect 32508 7588 32564 7756
rect 34850 7644 34860 7700
rect 34916 7644 36092 7700
rect 36148 7644 42028 7700
rect 42084 7644 42094 7700
rect 14550 7532 14588 7588
rect 14644 7532 14654 7588
rect 17602 7532 17612 7588
rect 17668 7532 19516 7588
rect 19572 7532 19582 7588
rect 19954 7532 19964 7588
rect 20020 7532 20692 7588
rect 25302 7532 25340 7588
rect 25396 7532 25406 7588
rect 26002 7532 26012 7588
rect 26068 7532 31948 7588
rect 32004 7532 32014 7588
rect 32498 7532 32508 7588
rect 32564 7532 32574 7588
rect 33506 7532 33516 7588
rect 33572 7532 34412 7588
rect 34468 7532 34478 7588
rect 10994 7420 11004 7476
rect 11060 7420 11676 7476
rect 11732 7420 13468 7476
rect 13524 7420 13534 7476
rect 15092 7420 15484 7476
rect 15540 7420 16156 7476
rect 16212 7420 16222 7476
rect 17938 7420 17948 7476
rect 18004 7420 18620 7476
rect 18676 7420 18686 7476
rect 20290 7420 20300 7476
rect 20356 7420 21644 7476
rect 21700 7420 21710 7476
rect 24098 7420 24108 7476
rect 24164 7420 26236 7476
rect 26292 7420 26302 7476
rect 27570 7420 27580 7476
rect 27636 7420 29708 7476
rect 29764 7420 29774 7476
rect 38994 7420 39004 7476
rect 39060 7420 42252 7476
rect 42308 7420 42318 7476
rect 49074 7420 49084 7476
rect 49140 7420 50876 7476
rect 50932 7420 50942 7476
rect 15092 7364 15148 7420
rect 13570 7308 13580 7364
rect 13636 7308 15148 7364
rect 16258 7308 16268 7364
rect 16324 7308 18508 7364
rect 18564 7308 18574 7364
rect 19394 7308 19404 7364
rect 19460 7308 23996 7364
rect 24052 7308 24062 7364
rect 24210 7308 24220 7364
rect 24276 7308 24286 7364
rect 24658 7308 24668 7364
rect 24724 7308 26012 7364
rect 26068 7308 26078 7364
rect 28018 7308 28028 7364
rect 28084 7308 41244 7364
rect 41300 7308 41310 7364
rect 47058 7308 47068 7364
rect 47124 7308 48300 7364
rect 48356 7308 49420 7364
rect 49476 7308 49486 7364
rect 24220 7252 24276 7308
rect 18722 7196 18732 7252
rect 18788 7196 19292 7252
rect 19348 7196 21980 7252
rect 22036 7196 22046 7252
rect 23874 7196 23884 7252
rect 23940 7196 24276 7252
rect 24546 7196 24556 7252
rect 24612 7196 24892 7252
rect 24948 7196 24958 7252
rect 25890 7084 25900 7140
rect 25956 7084 26124 7140
rect 26180 7084 26190 7140
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 10882 6972 10892 7028
rect 10948 6972 12236 7028
rect 12292 6972 12302 7028
rect 19282 6972 19292 7028
rect 19348 6972 19628 7028
rect 19684 6972 19694 7028
rect 21746 6972 21756 7028
rect 21812 6972 22204 7028
rect 22260 6972 22270 7028
rect 24882 6972 24892 7028
rect 24948 6972 25340 7028
rect 25396 6972 25406 7028
rect 25666 6972 25676 7028
rect 25732 6972 27244 7028
rect 27300 6972 27310 7028
rect 13990 6860 14028 6916
rect 14084 6860 14094 6916
rect 20850 6860 20860 6916
rect 20916 6860 26572 6916
rect 26628 6860 26638 6916
rect 9874 6748 9884 6804
rect 9940 6748 13468 6804
rect 13524 6748 13534 6804
rect 14466 6748 14476 6804
rect 14532 6748 18060 6804
rect 18116 6748 18126 6804
rect 18274 6748 18284 6804
rect 18340 6748 20748 6804
rect 20804 6748 21196 6804
rect 21252 6748 21262 6804
rect 24070 6748 24108 6804
rect 24164 6748 24174 6804
rect 24406 6748 24444 6804
rect 24500 6748 24510 6804
rect 28802 6748 28812 6804
rect 28868 6748 29260 6804
rect 29316 6748 29326 6804
rect 29810 6748 29820 6804
rect 29876 6748 32620 6804
rect 32676 6748 35644 6804
rect 35700 6748 35710 6804
rect 11890 6636 11900 6692
rect 11956 6636 13692 6692
rect 13748 6636 16044 6692
rect 16100 6636 16110 6692
rect 18386 6636 18396 6692
rect 18452 6636 20524 6692
rect 20580 6636 20590 6692
rect 21410 6636 21420 6692
rect 21476 6636 22092 6692
rect 22148 6636 22428 6692
rect 22484 6636 22494 6692
rect 26450 6636 26460 6692
rect 26516 6636 28476 6692
rect 28532 6636 31612 6692
rect 31668 6636 31678 6692
rect 32946 6636 32956 6692
rect 33012 6636 33964 6692
rect 34020 6636 34030 6692
rect 35858 6636 35868 6692
rect 35924 6636 38108 6692
rect 38164 6636 38174 6692
rect 38612 6580 38668 6692
rect 38724 6636 38734 6692
rect 11330 6524 11340 6580
rect 11396 6524 14700 6580
rect 14756 6524 15036 6580
rect 15092 6524 15708 6580
rect 15764 6524 15774 6580
rect 16482 6524 16492 6580
rect 16548 6524 18732 6580
rect 18788 6524 18798 6580
rect 19058 6524 19068 6580
rect 19124 6524 19852 6580
rect 19908 6524 21644 6580
rect 21700 6524 21710 6580
rect 24098 6524 24108 6580
rect 24164 6524 24444 6580
rect 24500 6524 24510 6580
rect 26226 6524 26236 6580
rect 26292 6524 28140 6580
rect 28196 6524 28206 6580
rect 28354 6524 28364 6580
rect 28420 6524 32508 6580
rect 32564 6524 32574 6580
rect 37426 6524 37436 6580
rect 37492 6524 38668 6580
rect 12674 6412 12684 6468
rect 12740 6412 15820 6468
rect 15876 6412 15886 6468
rect 18498 6412 18508 6468
rect 18564 6412 20468 6468
rect 20626 6412 20636 6468
rect 20692 6412 22428 6468
rect 22484 6412 22494 6468
rect 23762 6412 23772 6468
rect 23828 6412 24668 6468
rect 24724 6412 24734 6468
rect 26786 6412 26796 6468
rect 26852 6412 28812 6468
rect 28868 6412 28878 6468
rect 37314 6412 37324 6468
rect 37380 6412 38444 6468
rect 38500 6412 38510 6468
rect 20412 6356 20468 6412
rect 20412 6300 21084 6356
rect 21140 6300 21150 6356
rect 23650 6300 23660 6356
rect 23716 6300 25788 6356
rect 25844 6300 26348 6356
rect 26404 6300 26414 6356
rect 32162 6300 32172 6356
rect 32228 6300 35196 6356
rect 35252 6300 41468 6356
rect 41524 6300 41534 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 25330 6188 25340 6244
rect 25396 6188 26236 6244
rect 26292 6188 26302 6244
rect 12338 6076 12348 6132
rect 12404 6076 14476 6132
rect 14532 6076 14542 6132
rect 16930 6076 16940 6132
rect 16996 6076 17836 6132
rect 17892 6076 18956 6132
rect 19012 6076 19022 6132
rect 20178 6076 20188 6132
rect 20244 6076 27468 6132
rect 27524 6076 27534 6132
rect 29922 6076 29932 6132
rect 29988 6076 30604 6132
rect 30660 6076 30670 6132
rect 42802 6076 42812 6132
rect 42868 6076 44268 6132
rect 44324 6076 44334 6132
rect 15138 5964 15148 6020
rect 15204 5964 19852 6020
rect 19908 5964 19918 6020
rect 22614 5964 22652 6020
rect 22708 5964 22718 6020
rect 24322 5964 24332 6020
rect 24388 5964 24780 6020
rect 24836 5964 26684 6020
rect 26740 5964 26750 6020
rect 26898 5964 26908 6020
rect 26964 5964 27692 6020
rect 27748 5964 29036 6020
rect 29092 5964 29102 6020
rect 48738 5964 48748 6020
rect 48804 5964 49420 6020
rect 49476 5964 49486 6020
rect 15586 5852 15596 5908
rect 15652 5852 16268 5908
rect 16324 5852 16334 5908
rect 17266 5852 17276 5908
rect 17332 5852 18508 5908
rect 18564 5852 18574 5908
rect 19506 5852 19516 5908
rect 19572 5852 20412 5908
rect 20468 5852 20478 5908
rect 21634 5852 21644 5908
rect 21700 5852 22316 5908
rect 22372 5852 22382 5908
rect 22978 5852 22988 5908
rect 23044 5852 23772 5908
rect 23828 5852 23838 5908
rect 25890 5852 25900 5908
rect 25956 5852 25966 5908
rect 28130 5852 28140 5908
rect 28196 5852 29372 5908
rect 29428 5852 29438 5908
rect 36194 5852 36204 5908
rect 36260 5852 36876 5908
rect 36932 5852 36942 5908
rect 38434 5852 38444 5908
rect 38500 5852 39676 5908
rect 39732 5852 39742 5908
rect 40002 5852 40012 5908
rect 40068 5852 40348 5908
rect 40404 5852 41244 5908
rect 41300 5852 41310 5908
rect 43138 5852 43148 5908
rect 43204 5852 44604 5908
rect 44660 5852 44670 5908
rect 46050 5852 46060 5908
rect 46116 5852 46732 5908
rect 46788 5852 47628 5908
rect 47684 5852 47694 5908
rect 48402 5852 48412 5908
rect 48468 5852 48860 5908
rect 48916 5852 49644 5908
rect 49700 5852 49710 5908
rect 25900 5796 25956 5852
rect 44604 5796 44660 5852
rect 48412 5796 48468 5852
rect 16594 5740 16604 5796
rect 16660 5740 18060 5796
rect 18116 5740 20524 5796
rect 20580 5740 20590 5796
rect 21522 5740 21532 5796
rect 21588 5740 25956 5796
rect 37650 5740 37660 5796
rect 37716 5740 39452 5796
rect 39508 5740 39518 5796
rect 44604 5740 46508 5796
rect 46564 5740 46574 5796
rect 47282 5740 47292 5796
rect 47348 5740 48468 5796
rect 13122 5628 13132 5684
rect 13188 5628 14588 5684
rect 14644 5628 17276 5684
rect 17332 5628 17342 5684
rect 19282 5628 19292 5684
rect 19348 5628 19852 5684
rect 19908 5628 20860 5684
rect 20916 5628 20926 5684
rect 21298 5628 21308 5684
rect 21364 5628 23100 5684
rect 23156 5628 23166 5684
rect 42130 5628 42140 5684
rect 42196 5628 42924 5684
rect 42980 5628 42990 5684
rect 43698 5628 43708 5684
rect 43764 5628 44380 5684
rect 44436 5628 44446 5684
rect 48178 5628 48188 5684
rect 48244 5628 50092 5684
rect 50148 5628 50158 5684
rect 11890 5516 11900 5572
rect 11956 5516 12572 5572
rect 12628 5516 13468 5572
rect 13524 5516 15708 5572
rect 15764 5516 17388 5572
rect 17444 5516 17454 5572
rect 20290 5516 20300 5572
rect 20356 5516 21084 5572
rect 21140 5516 21150 5572
rect 24770 5516 24780 5572
rect 24836 5516 25340 5572
rect 25396 5516 25406 5572
rect 26898 5516 26908 5572
rect 26964 5516 29204 5572
rect 39778 5516 39788 5572
rect 39844 5516 40572 5572
rect 40628 5516 41468 5572
rect 41524 5516 41534 5572
rect 41906 5516 41916 5572
rect 41972 5516 46396 5572
rect 46452 5516 47852 5572
rect 47908 5516 47918 5572
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 14812 5404 16604 5460
rect 16660 5404 16670 5460
rect 16818 5404 16828 5460
rect 16884 5404 20524 5460
rect 20580 5404 21364 5460
rect 24098 5404 24108 5460
rect 24164 5404 28476 5460
rect 28532 5404 28542 5460
rect 14812 5348 14868 5404
rect 21308 5348 21364 5404
rect 12786 5292 12796 5348
rect 12852 5292 14812 5348
rect 14868 5292 14878 5348
rect 16380 5292 18284 5348
rect 18340 5292 18350 5348
rect 19730 5292 19740 5348
rect 19796 5292 20748 5348
rect 20804 5292 20814 5348
rect 21308 5292 24332 5348
rect 24388 5292 25228 5348
rect 25284 5292 25294 5348
rect 25442 5292 25452 5348
rect 25508 5292 25518 5348
rect 25778 5292 25788 5348
rect 25844 5292 27804 5348
rect 27860 5292 27870 5348
rect 28130 5292 28140 5348
rect 28196 5292 28812 5348
rect 28868 5292 28878 5348
rect 16380 5236 16436 5292
rect 25452 5236 25508 5292
rect 29148 5236 29204 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 40002 5404 40012 5460
rect 40068 5404 42364 5460
rect 42420 5404 42430 5460
rect 39442 5292 39452 5348
rect 39508 5292 40796 5348
rect 40852 5292 40862 5348
rect 14018 5180 14028 5236
rect 14084 5180 16436 5236
rect 18386 5180 18396 5236
rect 18452 5180 19516 5236
rect 19572 5180 20076 5236
rect 20132 5180 20142 5236
rect 20626 5180 20636 5236
rect 20692 5180 20972 5236
rect 21028 5180 21038 5236
rect 25452 5180 27020 5236
rect 27076 5180 27086 5236
rect 29138 5180 29148 5236
rect 29204 5180 29214 5236
rect 30370 5180 30380 5236
rect 30436 5180 31612 5236
rect 31668 5180 32732 5236
rect 32788 5180 32798 5236
rect 39106 5180 39116 5236
rect 39172 5180 42140 5236
rect 42196 5180 42206 5236
rect 44370 5180 44380 5236
rect 44436 5180 46732 5236
rect 46788 5180 48076 5236
rect 48132 5180 48142 5236
rect 15250 5068 15260 5124
rect 15316 5068 16604 5124
rect 16660 5068 17836 5124
rect 17892 5068 17902 5124
rect 18610 5068 18620 5124
rect 18676 5068 22204 5124
rect 22260 5068 22270 5124
rect 23202 5068 23212 5124
rect 23268 5068 25116 5124
rect 25172 5068 28140 5124
rect 28196 5068 28206 5124
rect 28466 5068 28476 5124
rect 28532 5068 29484 5124
rect 29540 5068 29550 5124
rect 38658 5068 38668 5124
rect 38724 5068 39004 5124
rect 39060 5068 39340 5124
rect 39396 5068 39406 5124
rect 40450 5068 40460 5124
rect 40516 5068 45164 5124
rect 45220 5068 45230 5124
rect 46050 5068 46060 5124
rect 46116 5068 47068 5124
rect 47124 5068 47134 5124
rect 50082 5068 50092 5124
rect 50148 5068 51212 5124
rect 51268 5068 51278 5124
rect 14018 4956 14028 5012
rect 14084 4956 14364 5012
rect 14420 4956 14430 5012
rect 18722 4956 18732 5012
rect 18788 4956 25452 5012
rect 25508 4956 25518 5012
rect 28130 4956 28140 5012
rect 28196 4956 29708 5012
rect 29764 4956 29774 5012
rect 34290 4956 34300 5012
rect 34356 4956 35644 5012
rect 35700 4956 35710 5012
rect 42130 4956 42140 5012
rect 42196 4956 43036 5012
rect 43092 4956 44044 5012
rect 44100 4956 44110 5012
rect 48962 4956 48972 5012
rect 49028 4956 51324 5012
rect 51380 4956 51390 5012
rect 14914 4844 14924 4900
rect 14980 4844 15820 4900
rect 15876 4844 15886 4900
rect 16370 4844 16380 4900
rect 16436 4844 16940 4900
rect 16996 4844 17006 4900
rect 17266 4844 17276 4900
rect 17332 4844 19292 4900
rect 19348 4844 19358 4900
rect 19506 4844 19516 4900
rect 19572 4844 20188 4900
rect 20244 4844 20254 4900
rect 22754 4844 22764 4900
rect 22820 4844 32116 4900
rect 32274 4844 32284 4900
rect 32340 4844 41916 4900
rect 41972 4844 41982 4900
rect 43652 4844 44156 4900
rect 44212 4844 45388 4900
rect 45444 4844 45454 4900
rect 50754 4844 50764 4900
rect 50820 4844 51436 4900
rect 51492 4844 51502 4900
rect 32060 4788 32116 4844
rect 14690 4732 14700 4788
rect 14756 4732 19684 4788
rect 22866 4732 22876 4788
rect 22932 4732 28140 4788
rect 28196 4732 28206 4788
rect 32060 4732 37884 4788
rect 37940 4732 37950 4788
rect 15250 4620 15260 4676
rect 15316 4620 19180 4676
rect 19236 4620 19246 4676
rect 17602 4508 17612 4564
rect 17668 4508 18060 4564
rect 18116 4508 18126 4564
rect 18386 4508 18396 4564
rect 18452 4508 19404 4564
rect 19460 4508 19470 4564
rect 18274 4396 18284 4452
rect 18340 4396 18844 4452
rect 18900 4396 18910 4452
rect 19254 4396 19292 4452
rect 19348 4396 19358 4452
rect 19628 4340 19684 4732
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 22754 4620 22764 4676
rect 22820 4620 25340 4676
rect 25396 4620 25406 4676
rect 30706 4620 30716 4676
rect 30772 4620 40460 4676
rect 40516 4620 40526 4676
rect 19954 4508 19964 4564
rect 20020 4508 21420 4564
rect 21476 4508 21486 4564
rect 21858 4508 21868 4564
rect 21924 4508 23324 4564
rect 23380 4508 23390 4564
rect 24322 4508 24332 4564
rect 24388 4508 25452 4564
rect 25508 4508 25518 4564
rect 30370 4508 30380 4564
rect 30436 4508 33068 4564
rect 33124 4508 33134 4564
rect 34066 4508 34076 4564
rect 34132 4508 35084 4564
rect 35140 4508 35532 4564
rect 35588 4508 35598 4564
rect 38434 4508 38444 4564
rect 38500 4508 39564 4564
rect 39620 4508 39630 4564
rect 43652 4452 43708 4844
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 45266 4620 45276 4676
rect 45332 4620 47404 4676
rect 47460 4620 49084 4676
rect 49140 4620 49644 4676
rect 49700 4620 49710 4676
rect 21522 4396 21532 4452
rect 21588 4396 22204 4452
rect 22260 4396 22876 4452
rect 22932 4396 22942 4452
rect 24434 4396 24444 4452
rect 24500 4396 25228 4452
rect 25284 4396 25294 4452
rect 25554 4396 25564 4452
rect 25620 4396 25630 4452
rect 34514 4396 34524 4452
rect 34580 4396 35308 4452
rect 35364 4396 35374 4452
rect 38994 4396 39004 4452
rect 39060 4396 42812 4452
rect 42868 4396 43708 4452
rect 25564 4340 25620 4396
rect 18582 4284 18620 4340
rect 18676 4284 18686 4340
rect 19628 4284 25620 4340
rect 30594 4284 30604 4340
rect 30660 4284 31836 4340
rect 31892 4284 31902 4340
rect 34290 4284 34300 4340
rect 34356 4284 34972 4340
rect 35028 4284 35038 4340
rect 15810 4172 15820 4228
rect 15876 4172 24444 4228
rect 24500 4172 24510 4228
rect 34402 4172 34412 4228
rect 34468 4172 38108 4228
rect 38164 4172 38174 4228
rect 19394 4060 19404 4116
rect 19460 4060 20524 4116
rect 20580 4060 20590 4116
rect 23090 4060 23100 4116
rect 23156 4060 26348 4116
rect 26404 4060 26414 4116
rect 35858 4060 35868 4116
rect 35924 4060 38668 4116
rect 43698 4060 43708 4116
rect 43764 4060 44940 4116
rect 44996 4060 45006 4116
rect 51090 4060 51100 4116
rect 51156 4060 52332 4116
rect 52388 4060 52398 4116
rect 38612 4004 38668 4060
rect 16930 3948 16940 4004
rect 16996 3948 21532 4004
rect 21588 3948 21598 4004
rect 38612 3948 47180 4004
rect 47236 3948 48860 4004
rect 48916 3948 48926 4004
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 12002 3836 12012 3892
rect 12068 3836 14700 3892
rect 14756 3836 16492 3892
rect 16548 3836 19292 3892
rect 19348 3836 19358 3892
rect 14578 3612 14588 3668
rect 14644 3612 15820 3668
rect 15876 3612 15886 3668
rect 19142 3612 19180 3668
rect 19236 3612 19246 3668
rect 28774 3612 28812 3668
rect 28868 3612 28878 3668
rect 42354 3612 42364 3668
rect 42420 3612 44604 3668
rect 44660 3612 44670 3668
rect 50418 3612 50428 3668
rect 50484 3612 52220 3668
rect 52276 3612 52286 3668
rect 15820 3556 15876 3612
rect 15820 3500 21980 3556
rect 22036 3500 23100 3556
rect 23156 3500 23166 3556
rect 28914 3388 28924 3444
rect 28980 3388 30044 3444
rect 30100 3388 30110 3444
rect 46386 3388 46396 3444
rect 46452 3388 48972 3444
rect 49028 3388 49038 3444
rect 4722 3276 4732 3332
rect 4788 3276 5516 3332
rect 5572 3276 5582 3332
rect 11554 3276 11564 3332
rect 11620 3276 19740 3332
rect 19796 3276 19806 3332
rect 20402 3276 20412 3332
rect 20468 3276 41132 3332
rect 41188 3276 41198 3332
rect 52434 3276 52444 3332
rect 52500 3276 54124 3332
rect 54180 3276 54190 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
rect 11890 2828 11900 2884
rect 11956 2828 25004 2884
rect 25060 2828 25070 2884
rect 13234 2716 13244 2772
rect 13300 2716 29148 2772
rect 29204 2716 29214 2772
rect 16594 2604 16604 2660
rect 16660 2604 27132 2660
rect 27188 2604 27198 2660
rect 15250 1596 15260 1652
rect 15316 1596 30492 1652
rect 30548 1596 30558 1652
rect 16706 1484 16716 1540
rect 16772 1484 27692 1540
rect 27748 1484 27758 1540
rect 14466 1372 14476 1428
rect 14532 1372 23884 1428
rect 23940 1372 23950 1428
<< via3 >>
rect 20524 57820 20580 57876
rect 12012 57596 12068 57652
rect 21420 56700 21476 56756
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 17836 55580 17892 55636
rect 15036 55244 15092 55300
rect 31724 55020 31780 55076
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 17836 54460 17892 54516
rect 15036 54348 15092 54404
rect 16268 54348 16324 54404
rect 30604 54348 30660 54404
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 15932 54012 15988 54068
rect 29820 53900 29876 53956
rect 23660 53676 23716 53732
rect 13356 53564 13412 53620
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 17612 53116 17668 53172
rect 33628 53116 33684 53172
rect 13356 53004 13412 53060
rect 13804 52780 13860 52836
rect 11788 52668 11844 52724
rect 23660 52668 23716 52724
rect 34524 52668 34580 52724
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 20748 52444 20804 52500
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 19068 52332 19124 52388
rect 14364 52220 14420 52276
rect 19628 52220 19684 52276
rect 20188 52220 20244 52276
rect 15484 51996 15540 52052
rect 30828 52108 30884 52164
rect 20636 51884 20692 51940
rect 20860 51884 20916 51940
rect 29260 51884 29316 51940
rect 31388 51884 31444 51940
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 18732 51324 18788 51380
rect 20300 51324 20356 51380
rect 20748 51324 20804 51380
rect 22876 51324 22932 51380
rect 24668 51324 24724 51380
rect 27132 51324 27188 51380
rect 31388 51100 31444 51156
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 20188 50876 20244 50932
rect 26684 50876 26740 50932
rect 24332 50540 24388 50596
rect 30044 50540 30100 50596
rect 30604 50428 30660 50484
rect 31388 50428 31444 50484
rect 20860 50204 20916 50260
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 18844 50092 18900 50148
rect 27244 49756 27300 49812
rect 27804 49644 27860 49700
rect 30828 49420 30884 49476
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 27580 49196 27636 49252
rect 20524 49084 20580 49140
rect 28364 48972 28420 49028
rect 19628 48860 19684 48916
rect 20300 48636 20356 48692
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 27804 48524 27860 48580
rect 27244 48412 27300 48468
rect 29820 48412 29876 48468
rect 27692 48188 27748 48244
rect 34524 48188 34580 48244
rect 18732 47964 18788 48020
rect 21420 47964 21476 48020
rect 27580 47964 27636 48020
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 26684 47740 26740 47796
rect 28364 47628 28420 47684
rect 29708 47628 29764 47684
rect 11788 47516 11844 47572
rect 29708 47292 29764 47348
rect 28476 47180 28532 47236
rect 18844 47068 18900 47124
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 19516 46956 19572 47012
rect 27244 46956 27300 47012
rect 24220 46844 24276 46900
rect 20524 46732 20580 46788
rect 27132 46732 27188 46788
rect 12012 46620 12068 46676
rect 26460 46620 26516 46676
rect 26684 46620 26740 46676
rect 27244 46620 27300 46676
rect 28476 46620 28532 46676
rect 6860 46508 6916 46564
rect 29596 46396 29652 46452
rect 29484 46284 29540 46340
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 28588 46060 28644 46116
rect 18732 45948 18788 46004
rect 23884 45948 23940 46004
rect 29932 45948 29988 46004
rect 34300 45836 34356 45892
rect 29148 45724 29204 45780
rect 13804 45500 13860 45556
rect 17388 45500 17444 45556
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 14812 45388 14868 45444
rect 19180 45388 19236 45444
rect 21532 45276 21588 45332
rect 19516 45164 19572 45220
rect 25900 44940 25956 44996
rect 13804 44828 13860 44884
rect 15484 44828 15540 44884
rect 34188 44828 34244 44884
rect 29036 44716 29092 44772
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 24556 44492 24612 44548
rect 28700 44492 28756 44548
rect 29260 44492 29316 44548
rect 18956 44268 19012 44324
rect 26460 44268 26516 44324
rect 19628 44156 19684 44212
rect 20524 44156 20580 44212
rect 14476 44044 14532 44100
rect 23100 44044 23156 44100
rect 26012 44044 26068 44100
rect 29484 44268 29540 44324
rect 27020 44044 27076 44100
rect 34188 43932 34244 43988
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 20636 43708 20692 43764
rect 29260 43708 29316 43764
rect 34972 43708 35028 43764
rect 22316 43596 22372 43652
rect 22876 43596 22932 43652
rect 25788 43596 25844 43652
rect 29036 43484 29092 43540
rect 28700 43372 28756 43428
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 16268 42924 16324 42980
rect 27356 42924 27412 42980
rect 30044 42924 30100 42980
rect 18732 42700 18788 42756
rect 26796 42700 26852 42756
rect 27356 42700 27412 42756
rect 30716 42476 30772 42532
rect 26796 42364 26852 42420
rect 46508 42364 46564 42420
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 22204 42140 22260 42196
rect 24332 42140 24388 42196
rect 26684 42140 26740 42196
rect 23660 42028 23716 42084
rect 14588 41916 14644 41972
rect 17388 41916 17444 41972
rect 29596 41916 29652 41972
rect 46508 41580 46564 41636
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 23436 41468 23492 41524
rect 25228 41132 25284 41188
rect 28588 41132 28644 41188
rect 29708 41132 29764 41188
rect 24220 41020 24276 41076
rect 25676 40908 25732 40964
rect 13356 40796 13412 40852
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 12012 40572 12068 40628
rect 22204 40572 22260 40628
rect 33068 40572 33124 40628
rect 19180 40348 19236 40404
rect 24668 40236 24724 40292
rect 14364 40012 14420 40068
rect 14700 40012 14756 40068
rect 33852 40012 33908 40068
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 29484 39788 29540 39844
rect 23884 39676 23940 39732
rect 25676 39452 25732 39508
rect 18956 39340 19012 39396
rect 14700 39228 14756 39284
rect 19516 39228 19572 39284
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 23884 39340 23940 39396
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 33852 39116 33908 39172
rect 33628 39004 33684 39060
rect 11788 38668 11844 38724
rect 14588 38668 14644 38724
rect 19516 38668 19572 38724
rect 23100 38668 23156 38724
rect 29260 38556 29316 38612
rect 19180 38444 19236 38500
rect 21532 38444 21588 38500
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 25228 38332 25284 38388
rect 11788 38220 11844 38276
rect 25900 38220 25956 38276
rect 22316 38108 22372 38164
rect 27692 38108 27748 38164
rect 18732 37996 18788 38052
rect 29484 37996 29540 38052
rect 33068 37996 33124 38052
rect 19628 37884 19684 37940
rect 26012 37772 26068 37828
rect 27020 37660 27076 37716
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 15932 37436 15988 37492
rect 17612 37436 17668 37492
rect 26460 37212 26516 37268
rect 24556 36876 24612 36932
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 29148 36764 29204 36820
rect 34300 36652 34356 36708
rect 14476 36428 14532 36484
rect 26460 36428 26516 36484
rect 30716 36316 30772 36372
rect 19516 36092 19572 36148
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 23436 35980 23492 36036
rect 34972 35980 35028 36036
rect 14476 35868 14532 35924
rect 25788 35756 25844 35812
rect 6860 35532 6916 35588
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 15036 35196 15092 35252
rect 14812 35084 14868 35140
rect 29932 34524 29988 34580
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 19068 34412 19124 34468
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19068 32956 19124 33012
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 19180 32844 19236 32900
rect 31724 32732 31780 32788
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 31388 31836 31444 31892
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 26572 30828 26628 30884
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 28700 30492 28756 30548
rect 11676 30268 11732 30324
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 27580 29484 27636 29540
rect 16716 29260 16772 29316
rect 18732 29148 18788 29204
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 11004 28924 11060 28980
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 20636 28252 20692 28308
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 16268 28028 16324 28084
rect 16940 27916 16996 27972
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 18508 27132 18564 27188
rect 28812 26908 28868 26964
rect 19404 26684 19460 26740
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 19404 26460 19460 26516
rect 14364 26124 14420 26180
rect 16380 26124 16436 26180
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 14364 25788 14420 25844
rect 31836 25228 31892 25284
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 16716 24780 16772 24836
rect 28700 24780 28756 24836
rect 23772 24556 23828 24612
rect 11004 24444 11060 24500
rect 18732 24332 18788 24388
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19404 23772 19460 23828
rect 20412 23772 20468 23828
rect 31612 23772 31668 23828
rect 11228 23660 11284 23716
rect 16828 23660 16884 23716
rect 22428 23660 22484 23716
rect 31612 23548 31668 23604
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 26460 23324 26516 23380
rect 16268 23100 16324 23156
rect 15596 22988 15652 23044
rect 26012 22764 26068 22820
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 18508 22540 18564 22596
rect 17836 22428 17892 22484
rect 23436 22316 23492 22372
rect 26684 22316 26740 22372
rect 13916 22204 13972 22260
rect 16380 22204 16436 22260
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 17836 21868 17892 21924
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 26460 21756 26516 21812
rect 14364 21644 14420 21700
rect 26012 21644 26068 21700
rect 23884 21420 23940 21476
rect 7868 21196 7924 21252
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 26684 21084 26740 21140
rect 20636 20748 20692 20804
rect 31948 20636 32004 20692
rect 24556 20524 24612 20580
rect 19292 20412 19348 20468
rect 25004 20412 25060 20468
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 31948 20412 32004 20468
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 11900 20300 11956 20356
rect 16268 20300 16324 20356
rect 12684 20188 12740 20244
rect 11676 20076 11732 20132
rect 15372 20076 15428 20132
rect 11676 19852 11732 19908
rect 17500 19852 17556 19908
rect 18172 19740 18228 19796
rect 14364 19628 14420 19684
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 10668 19404 10724 19460
rect 18172 19404 18228 19460
rect 21980 19292 22036 19348
rect 9324 19180 9380 19236
rect 26012 19180 26068 19236
rect 17052 19068 17108 19124
rect 22652 19068 22708 19124
rect 23548 19068 23604 19124
rect 9548 18956 9604 19012
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 7756 18620 7812 18676
rect 16380 18508 16436 18564
rect 16716 18508 16772 18564
rect 9324 18396 9380 18452
rect 17388 18396 17444 18452
rect 23436 18396 23492 18452
rect 12684 18284 12740 18340
rect 10668 18172 10724 18228
rect 19628 18172 19684 18228
rect 27692 18284 27748 18340
rect 19516 18060 19572 18116
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 23324 17836 23380 17892
rect 11004 17612 11060 17668
rect 14476 17388 14532 17444
rect 24556 17276 24612 17332
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 13916 17164 13972 17220
rect 23996 17052 24052 17108
rect 8428 16940 8484 16996
rect 24668 16940 24724 16996
rect 20860 16828 20916 16884
rect 11228 16604 11284 16660
rect 11900 16604 11956 16660
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 17500 16380 17556 16436
rect 20636 16380 20692 16436
rect 25116 16380 25172 16436
rect 26684 16268 26740 16324
rect 11340 16156 11396 16212
rect 19292 16156 19348 16212
rect 17612 15820 17668 15876
rect 22988 15820 23044 15876
rect 23996 15820 24052 15876
rect 21980 15708 22036 15764
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 15036 15596 15092 15652
rect 31500 15596 31556 15652
rect 11788 15484 11844 15540
rect 24668 15484 24724 15540
rect 9324 15372 9380 15428
rect 15092 15372 15148 15428
rect 17052 15372 17108 15428
rect 17388 15372 17444 15428
rect 21420 15372 21476 15428
rect 26012 15372 26068 15428
rect 22764 15260 22820 15316
rect 9548 15148 9604 15204
rect 11900 15148 11956 15204
rect 22428 15148 22484 15204
rect 15260 15036 15316 15092
rect 20188 15036 20244 15092
rect 8428 14924 8484 14980
rect 23660 14924 23716 14980
rect 28140 14924 28196 14980
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19628 14812 19684 14868
rect 12684 14588 12740 14644
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 24220 14140 24276 14196
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 23996 14028 24052 14084
rect 7756 13916 7812 13972
rect 23324 13916 23380 13972
rect 23548 13916 23604 13972
rect 16828 13804 16884 13860
rect 23660 13804 23716 13860
rect 11340 13692 11396 13748
rect 18396 13692 18452 13748
rect 20860 13692 20916 13748
rect 15372 13580 15428 13636
rect 16380 13468 16436 13524
rect 18060 13468 18116 13524
rect 21420 13468 21476 13524
rect 26684 13468 26740 13524
rect 7868 13356 7924 13412
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 22764 13244 22820 13300
rect 18396 13132 18452 13188
rect 25116 13132 25172 13188
rect 24220 13020 24276 13076
rect 22428 12908 22484 12964
rect 17612 12796 17668 12852
rect 22876 12572 22932 12628
rect 31500 12572 31556 12628
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 28140 12460 28196 12516
rect 17836 12348 17892 12404
rect 16268 12124 16324 12180
rect 27356 12124 27412 12180
rect 27580 12124 27636 12180
rect 11788 12012 11844 12068
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 22876 11900 22932 11956
rect 13580 11788 13636 11844
rect 16940 11788 16996 11844
rect 21868 11788 21924 11844
rect 27356 11788 27412 11844
rect 36988 11788 37044 11844
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 13580 11564 13636 11620
rect 24332 11564 24388 11620
rect 18396 11452 18452 11508
rect 15036 11340 15092 11396
rect 24108 11340 24164 11396
rect 24556 11340 24612 11396
rect 19404 11116 19460 11172
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 24556 11116 24612 11172
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 22988 10780 23044 10836
rect 25340 10780 25396 10836
rect 15596 10668 15652 10724
rect 18060 10668 18116 10724
rect 19628 10668 19684 10724
rect 23772 10668 23828 10724
rect 25788 10668 25844 10724
rect 31836 10668 31892 10724
rect 26348 10556 26404 10612
rect 29148 10444 29204 10500
rect 18396 10220 18452 10276
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19292 10108 19348 10164
rect 11676 9996 11732 10052
rect 25004 9996 25060 10052
rect 36988 9996 37044 10052
rect 14700 9884 14756 9940
rect 19404 9548 19460 9604
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 24332 9324 24388 9380
rect 19180 9212 19236 9268
rect 26124 9212 26180 9268
rect 26572 9212 26628 9268
rect 24108 9100 24164 9156
rect 18620 8764 18676 8820
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19628 8428 19684 8484
rect 14924 8316 14980 8372
rect 43708 8316 43764 8372
rect 15036 8204 15092 8260
rect 43708 8092 43764 8148
rect 21868 7980 21924 8036
rect 26348 7980 26404 8036
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 20972 7756 21028 7812
rect 20412 7644 20468 7700
rect 25788 7644 25844 7700
rect 14588 7532 14644 7588
rect 19516 7532 19572 7588
rect 25340 7532 25396 7588
rect 26124 7084 26180 7140
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19292 6972 19348 7028
rect 14028 6860 14084 6916
rect 24108 6748 24164 6804
rect 24444 6748 24500 6804
rect 22428 6636 22484 6692
rect 15036 6524 15092 6580
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 22652 5964 22708 6020
rect 19292 5628 19348 5684
rect 25340 5516 25396 5572
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 28140 5292 28196 5348
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 20972 5180 21028 5236
rect 28140 5068 28196 5124
rect 14028 4956 14084 5012
rect 14700 4732 14756 4788
rect 18060 4508 18116 4564
rect 19404 4508 19460 4564
rect 19292 4396 19348 4452
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 24444 4396 24500 4452
rect 18620 4284 18676 4340
rect 24444 4172 24500 4228
rect 19404 4060 19460 4116
rect 26348 4060 26404 4116
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 14588 3612 14644 3668
rect 19180 3612 19236 3668
rect 28812 3612 28868 3668
rect 20412 3276 20468 3332
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
rect 29148 2716 29204 2772
rect 15260 1596 15316 1652
rect 16716 1484 16772 1540
rect 27692 1484 27748 1540
rect 14476 1372 14532 1428
rect 23884 1372 23940 1428
<< metal4 >>
rect 20524 57876 20580 57886
rect 12012 57652 12068 57662
rect 4448 55692 4768 56508
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 11788 52724 11844 52734
rect 11788 47572 11844 52668
rect 11788 47506 11844 47516
rect 12012 46676 12068 57596
rect 19808 56476 20128 56508
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 17836 55636 17892 55646
rect 15036 55300 15092 55310
rect 15036 54404 15092 55244
rect 17836 54516 17892 55580
rect 17836 54450 17892 54460
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 6860 46564 6916 46574
rect 6860 35588 6916 46508
rect 12012 40628 12068 46620
rect 13356 53620 13412 53630
rect 13356 53060 13412 53564
rect 13356 40852 13412 53004
rect 13804 52836 13860 52846
rect 13804 45556 13860 52780
rect 13804 44884 13860 45500
rect 13804 44818 13860 44828
rect 14364 52276 14420 52286
rect 13356 40786 13412 40796
rect 12012 40562 12068 40572
rect 14364 40068 14420 52220
rect 14812 45444 14868 45454
rect 14364 40002 14420 40012
rect 14476 44100 14532 44110
rect 11788 38724 11844 38734
rect 11788 38276 11844 38668
rect 11788 38210 11844 38220
rect 14476 36484 14532 44044
rect 14588 41972 14644 41982
rect 14588 38724 14644 41916
rect 14700 40068 14756 40078
rect 14700 39284 14756 40012
rect 14700 39218 14756 39228
rect 14588 38658 14644 38668
rect 14476 35924 14532 36428
rect 14476 35858 14532 35868
rect 6860 35522 6916 35532
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 14812 35140 14868 45388
rect 15036 35252 15092 54348
rect 16268 54404 16324 54414
rect 15932 54068 15988 54078
rect 15484 52052 15540 52062
rect 15484 44884 15540 51996
rect 15484 44818 15540 44828
rect 15932 37492 15988 54012
rect 16268 42980 16324 54348
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 17612 53172 17668 53182
rect 16268 42914 16324 42924
rect 17388 45556 17444 45566
rect 17388 41972 17444 45500
rect 17388 41906 17444 41916
rect 15932 37426 15988 37436
rect 17612 37492 17668 53116
rect 19068 52388 19124 52398
rect 18732 51380 18788 51390
rect 18732 48020 18788 51324
rect 18732 47954 18788 47964
rect 18844 50148 18900 50158
rect 18844 47124 18900 50092
rect 18844 47058 18900 47068
rect 18732 46004 18788 46014
rect 18732 42756 18788 45948
rect 18732 38052 18788 42700
rect 18956 44324 19012 44334
rect 18956 39396 19012 44268
rect 18956 39330 19012 39340
rect 18732 37986 18788 37996
rect 17612 37426 17668 37436
rect 15036 35186 15092 35196
rect 14812 35074 14868 35084
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 19068 34468 19124 52332
rect 19628 52276 19684 52286
rect 19628 48916 19684 52220
rect 19628 48850 19684 48860
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 20188 52276 20244 52286
rect 20188 50932 20244 52220
rect 20188 50866 20244 50876
rect 20300 51380 20356 51390
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 20300 48692 20356 51324
rect 20524 49140 20580 57820
rect 21420 56756 21476 56766
rect 20748 52500 20804 52510
rect 20524 49074 20580 49084
rect 20636 51940 20692 51950
rect 20300 48626 20356 48636
rect 19808 47068 20128 48580
rect 19516 47012 19572 47022
rect 19180 45444 19236 45454
rect 19180 40404 19236 45388
rect 19180 40338 19236 40348
rect 19516 45220 19572 46956
rect 19516 39284 19572 45164
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19516 39218 19572 39228
rect 19628 44212 19684 44222
rect 19516 38724 19572 38734
rect 19068 33012 19124 34412
rect 19068 32946 19124 32956
rect 19180 38500 19236 38510
rect 19180 32900 19236 38444
rect 19516 36148 19572 38668
rect 19628 37940 19684 44156
rect 19628 37874 19684 37884
rect 19808 43932 20128 45444
rect 20524 46788 20580 46798
rect 20524 44212 20580 46732
rect 20524 44146 20580 44156
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19516 36082 19572 36092
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19180 32834 19236 32844
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 11676 30324 11732 30334
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 11004 28980 11060 28990
rect 11004 24500 11060 28924
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 7868 21252 7924 21262
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 7756 18676 7812 18686
rect 7756 13972 7812 18620
rect 7756 13906 7812 13916
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 7868 13412 7924 21196
rect 10668 19460 10724 19470
rect 9324 19236 9380 19246
rect 9324 18452 9380 19180
rect 8428 16996 8484 17006
rect 8428 14980 8484 16940
rect 9324 15428 9380 18396
rect 9324 15362 9380 15372
rect 9548 19012 9604 19022
rect 9548 15204 9604 18956
rect 10668 18228 10724 19404
rect 10668 18162 10724 18172
rect 11004 17668 11060 24444
rect 11004 17602 11060 17612
rect 11228 23716 11284 23726
rect 11228 16660 11284 23660
rect 11676 20132 11732 30268
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 16716 29316 16772 29326
rect 16268 28084 16324 28094
rect 14364 26180 14420 26190
rect 14364 25844 14420 26124
rect 14364 25778 14420 25788
rect 16268 23156 16324 28028
rect 16268 23090 16324 23100
rect 16380 26180 16436 26190
rect 15596 23044 15652 23054
rect 13916 22260 13972 22270
rect 11676 20066 11732 20076
rect 11900 20356 11956 20366
rect 11228 16594 11284 16604
rect 11676 19908 11732 19918
rect 9548 15138 9604 15148
rect 11340 16212 11396 16222
rect 8428 14914 8484 14924
rect 11340 13748 11396 16156
rect 11340 13682 11396 13692
rect 7868 13346 7924 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 11676 10052 11732 19852
rect 11900 16660 11956 20300
rect 11788 15540 11844 15550
rect 11788 12068 11844 15484
rect 11900 15204 11956 16604
rect 11900 15138 11956 15148
rect 12684 20244 12740 20254
rect 12684 18340 12740 20188
rect 12684 14644 12740 18284
rect 13916 17220 13972 22204
rect 14364 21700 14420 21710
rect 14364 19684 14420 21644
rect 14364 19618 14420 19628
rect 15372 20132 15428 20142
rect 13916 17154 13972 17164
rect 14476 17444 14532 17454
rect 12684 14578 12740 14588
rect 11788 12002 11844 12012
rect 13580 11844 13636 11854
rect 13580 11620 13636 11788
rect 13580 11554 13636 11564
rect 11676 9986 11732 9996
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 14028 6916 14084 6926
rect 14028 5012 14084 6860
rect 14028 4946 14084 4956
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 14476 1428 14532 17388
rect 15036 15652 15092 15662
rect 15036 15438 15092 15596
rect 15036 15428 15148 15438
rect 15036 15372 15092 15428
rect 15036 15362 15148 15372
rect 15036 11396 15092 15362
rect 14700 9940 14756 9950
rect 14588 7588 14644 7598
rect 14588 3668 14644 7532
rect 14700 4788 14756 9884
rect 15036 8398 15092 11340
rect 14924 8372 15092 8398
rect 14980 8342 15092 8372
rect 15260 15092 15316 15102
rect 14924 8306 14980 8316
rect 15036 8260 15092 8270
rect 15036 6580 15092 8204
rect 15036 6514 15092 6524
rect 14700 4722 14756 4732
rect 14588 3602 14644 3612
rect 15260 1652 15316 15036
rect 15372 13636 15428 20076
rect 15372 13570 15428 13580
rect 15596 10724 15652 22988
rect 16380 22260 16436 26124
rect 16716 24836 16772 29260
rect 18732 29204 18788 29214
rect 16716 24770 16772 24780
rect 16940 27972 16996 27982
rect 16268 20356 16324 20366
rect 16268 12180 16324 20300
rect 16380 18564 16436 22204
rect 16828 23716 16884 23726
rect 16380 13524 16436 18508
rect 16380 13458 16436 13468
rect 16716 18564 16772 18574
rect 16268 12114 16324 12124
rect 15596 10658 15652 10668
rect 15260 1586 15316 1596
rect 16716 1540 16772 18508
rect 16828 13860 16884 23660
rect 16828 13794 16884 13804
rect 16940 11844 16996 27916
rect 18508 27188 18564 27198
rect 18508 22596 18564 27132
rect 18732 24388 18788 29148
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 20636 43764 20692 51884
rect 20748 51380 20804 52444
rect 20748 51314 20804 51324
rect 20860 51940 20916 51950
rect 20860 50260 20916 51884
rect 20860 50194 20916 50204
rect 21420 48020 21476 56700
rect 35168 55692 35488 56508
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 31724 55076 31780 55086
rect 30604 54404 30660 54414
rect 29820 53956 29876 53966
rect 23660 53732 23716 53742
rect 23660 52724 23716 53676
rect 21420 47954 21476 47964
rect 22876 51380 22932 51390
rect 20636 28308 20692 43708
rect 21532 45332 21588 45342
rect 21532 38500 21588 45276
rect 22316 43652 22372 43662
rect 22204 42196 22260 42206
rect 22204 40628 22260 42140
rect 22204 40562 22260 40572
rect 21532 38434 21588 38444
rect 22316 38164 22372 43596
rect 22876 43652 22932 51324
rect 22876 43586 22932 43596
rect 23100 44100 23156 44110
rect 23100 38724 23156 44044
rect 23660 42084 23716 52668
rect 29260 51940 29316 51950
rect 24668 51380 24724 51390
rect 24332 50596 24388 50606
rect 24220 46900 24276 46910
rect 23660 42018 23716 42028
rect 23884 46004 23940 46014
rect 23100 38658 23156 38668
rect 23436 41524 23492 41534
rect 22316 38098 22372 38108
rect 23436 36036 23492 41468
rect 23884 39732 23940 45948
rect 24220 41076 24276 46844
rect 24332 42196 24388 50540
rect 24332 42130 24388 42140
rect 24556 44548 24612 44558
rect 24220 41010 24276 41020
rect 23884 39396 23940 39676
rect 23884 39330 23940 39340
rect 24556 36932 24612 44492
rect 24668 40292 24724 51324
rect 27132 51380 27188 51390
rect 26684 50932 26740 50942
rect 26684 47796 26740 50876
rect 26684 47730 26740 47740
rect 27132 46788 27188 51324
rect 27244 49812 27300 49822
rect 27244 48468 27300 49756
rect 27804 49700 27860 49710
rect 27244 48402 27300 48412
rect 27580 49252 27636 49262
rect 27580 48020 27636 49196
rect 27804 48580 27860 49644
rect 27804 48514 27860 48524
rect 28364 49028 28420 49038
rect 27580 47954 27636 47964
rect 27692 48244 27748 48254
rect 27132 46722 27188 46732
rect 27244 47012 27300 47022
rect 26460 46676 26516 46686
rect 25900 44996 25956 45006
rect 25788 43652 25844 43662
rect 24668 40226 24724 40236
rect 25228 41188 25284 41198
rect 25228 38388 25284 41132
rect 25676 40964 25732 40974
rect 25676 39508 25732 40908
rect 25676 39442 25732 39452
rect 25228 38322 25284 38332
rect 24556 36866 24612 36876
rect 23436 35970 23492 35980
rect 25788 35812 25844 43596
rect 25900 38276 25956 44940
rect 26460 44324 26516 46620
rect 25900 38210 25956 38220
rect 26012 44100 26068 44110
rect 26012 37828 26068 44044
rect 26012 37762 26068 37772
rect 26460 37268 26516 44268
rect 26684 46676 26740 46686
rect 26684 42196 26740 46620
rect 27244 46676 27300 46956
rect 27244 46610 27300 46620
rect 27020 44100 27076 44110
rect 26796 42756 26852 42766
rect 26796 42420 26852 42700
rect 26796 42354 26852 42364
rect 26684 42130 26740 42140
rect 27020 37716 27076 44044
rect 27356 42980 27412 42990
rect 27356 42756 27412 42924
rect 27356 42690 27412 42700
rect 27692 38164 27748 48188
rect 28364 47684 28420 48972
rect 28364 47618 28420 47628
rect 28476 47236 28532 47246
rect 28476 46676 28532 47180
rect 28476 46610 28532 46620
rect 28588 46116 28644 46126
rect 28588 41188 28644 46060
rect 29148 45780 29204 45790
rect 29036 44772 29092 44782
rect 28700 44548 28756 44558
rect 28700 43428 28756 44492
rect 29036 43540 29092 44716
rect 29036 43474 29092 43484
rect 28700 43362 28756 43372
rect 28588 41122 28644 41132
rect 27692 38098 27748 38108
rect 27020 37650 27076 37660
rect 26460 36484 26516 37212
rect 29148 36820 29204 45724
rect 29260 44548 29316 51884
rect 29820 48468 29876 53900
rect 29820 48402 29876 48412
rect 30044 50596 30100 50606
rect 29708 47684 29764 47694
rect 29708 47348 29764 47628
rect 29596 46452 29652 46462
rect 29260 44482 29316 44492
rect 29484 46340 29540 46350
rect 29484 44324 29540 46284
rect 29484 44258 29540 44268
rect 29260 43764 29316 43774
rect 29260 38612 29316 43708
rect 29596 41972 29652 46396
rect 29596 41906 29652 41916
rect 29708 41188 29764 47292
rect 29708 41122 29764 41132
rect 29932 46004 29988 46014
rect 29260 38546 29316 38556
rect 29484 39844 29540 39854
rect 29484 38052 29540 39788
rect 29484 37986 29540 37996
rect 29148 36754 29204 36764
rect 26460 36418 26516 36428
rect 25788 35746 25844 35756
rect 29932 34580 29988 45948
rect 30044 42980 30100 50540
rect 30604 50484 30660 54348
rect 30604 50418 30660 50428
rect 30828 52164 30884 52174
rect 30828 49476 30884 52108
rect 30828 49410 30884 49420
rect 31388 51940 31444 51950
rect 31388 51156 31444 51884
rect 31388 50484 31444 51100
rect 30044 42914 30100 42924
rect 30716 42532 30772 42542
rect 30716 36372 30772 42476
rect 30716 36306 30772 36316
rect 29932 34514 29988 34524
rect 31388 31892 31444 50428
rect 31724 32788 31780 55020
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 33628 53172 33684 53182
rect 33068 40628 33124 40638
rect 33068 38052 33124 40572
rect 33628 39060 33684 53116
rect 34524 52724 34580 52734
rect 34524 48244 34580 52668
rect 34524 48178 34580 48188
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 34300 45892 34356 45902
rect 34188 44884 34244 44894
rect 34188 43988 34244 44828
rect 34188 43922 34244 43932
rect 33852 40068 33908 40078
rect 33852 39172 33908 40012
rect 33852 39106 33908 39116
rect 33628 38994 33684 39004
rect 33068 37986 33124 37996
rect 34300 36708 34356 45836
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 34300 36642 34356 36652
rect 34972 43764 35028 43774
rect 34972 36036 35028 43708
rect 34972 35970 35028 35980
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 50528 56476 50848 56508
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 46508 42420 46564 42430
rect 46508 41636 46564 42364
rect 46508 41570 46564 41580
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 31724 32722 31780 32732
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 31388 31826 31444 31836
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 20636 28242 20692 28252
rect 26572 30884 26628 30894
rect 18732 24322 18788 24332
rect 19404 26740 19460 26750
rect 19404 26516 19460 26684
rect 19404 23828 19460 26460
rect 19404 23548 19460 23772
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 23772 24612 23828 24622
rect 19404 23492 19572 23548
rect 18508 22530 18564 22540
rect 17836 22484 17892 22494
rect 17836 21924 17892 22428
rect 17500 19908 17556 19918
rect 17052 19124 17108 19134
rect 17052 15428 17108 19068
rect 17052 15362 17108 15372
rect 17388 18452 17444 18462
rect 17388 15428 17444 18396
rect 17500 16436 17556 19852
rect 17500 16370 17556 16380
rect 17388 15362 17444 15372
rect 17612 15876 17668 15886
rect 17612 12852 17668 15820
rect 17612 12786 17668 12796
rect 17836 12404 17892 21868
rect 19292 20468 19348 20478
rect 18172 19796 18228 19806
rect 18172 19460 18228 19740
rect 18172 19394 18228 19404
rect 19292 16212 19348 20412
rect 19292 16146 19348 16156
rect 19516 18116 19572 23492
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 18396 13748 18452 13758
rect 17836 12338 17892 12348
rect 18060 13524 18116 13534
rect 16940 11778 16996 11788
rect 18060 10724 18116 13468
rect 18396 13188 18452 13692
rect 18396 13122 18452 13132
rect 18060 4564 18116 10668
rect 18396 11508 18452 11518
rect 18396 10276 18452 11452
rect 18396 10210 18452 10220
rect 19404 11172 19460 11182
rect 19292 10164 19348 10174
rect 19180 9268 19236 9278
rect 18060 4498 18116 4508
rect 18620 8820 18676 8830
rect 18620 4340 18676 8764
rect 18620 4274 18676 4284
rect 19180 3668 19236 9212
rect 19292 7028 19348 10108
rect 19292 6962 19348 6972
rect 19404 9604 19460 11116
rect 19292 5684 19348 5694
rect 19292 4452 19348 5628
rect 19292 4386 19348 4396
rect 19404 4564 19460 9548
rect 19516 7588 19572 18060
rect 19628 18228 19684 18238
rect 19628 14868 19684 18172
rect 19628 14802 19684 14812
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 20412 23828 20468 23838
rect 20412 17038 20468 23772
rect 22428 23716 22484 23726
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 20188 16982 20468 17038
rect 20636 20804 20692 20814
rect 20188 15092 20244 16982
rect 20636 16436 20692 20748
rect 21980 19348 22036 19358
rect 20636 16370 20692 16380
rect 20860 16884 20916 16894
rect 20188 15026 20244 15036
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 20860 13748 20916 16828
rect 21980 15764 22036 19292
rect 21980 15698 22036 15708
rect 20860 13682 20916 13692
rect 21420 15428 21476 15438
rect 21420 13524 21476 15372
rect 21420 13458 21476 13468
rect 22428 15204 22484 23660
rect 23436 22372 23492 22382
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 22428 12964 22484 15148
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19628 10724 19684 10734
rect 19628 8484 19684 10668
rect 19628 8418 19684 8428
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19516 7522 19572 7532
rect 19808 7868 20128 9380
rect 21868 11844 21924 11854
rect 21868 8036 21924 11788
rect 21868 7970 21924 7980
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19404 4116 19460 4508
rect 19404 4050 19460 4060
rect 19808 6300 20128 7812
rect 20972 7812 21028 7822
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19180 3602 19236 3612
rect 19808 3164 20128 4676
rect 20412 7700 20468 7710
rect 20412 3332 20468 7644
rect 20972 5236 21028 7756
rect 22428 6692 22484 12908
rect 22428 6626 22484 6636
rect 22652 19124 22708 19134
rect 22652 6020 22708 19068
rect 23436 18452 23492 22316
rect 23436 18386 23492 18396
rect 23548 19124 23604 19134
rect 23324 17892 23380 17902
rect 22988 15876 23044 15886
rect 22764 15316 22820 15326
rect 22764 13300 22820 15260
rect 22764 13234 22820 13244
rect 22876 12628 22932 12638
rect 22876 11956 22932 12572
rect 22876 11890 22932 11900
rect 22988 10836 23044 15820
rect 23324 13972 23380 17836
rect 23324 13906 23380 13916
rect 23548 13972 23604 19068
rect 23548 13906 23604 13916
rect 23660 14980 23716 14990
rect 23660 13860 23716 14924
rect 23660 13794 23716 13804
rect 22988 10770 23044 10780
rect 23772 10724 23828 24556
rect 26460 23380 26516 23390
rect 26012 22820 26068 22830
rect 26012 21700 26068 22764
rect 26460 21812 26516 23324
rect 26460 21746 26516 21756
rect 23772 10658 23828 10668
rect 23884 21476 23940 21486
rect 22652 5954 22708 5964
rect 20972 5170 21028 5180
rect 20412 3266 20468 3276
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 16716 1474 16772 1484
rect 14476 1362 14532 1372
rect 23884 1428 23940 21420
rect 24556 20580 24612 20590
rect 24556 17332 24612 20524
rect 24556 17266 24612 17276
rect 25004 20468 25060 20478
rect 23996 17108 24052 17118
rect 23996 15876 24052 17052
rect 23996 14084 24052 15820
rect 24668 16996 24724 17006
rect 24668 15540 24724 16940
rect 24668 15474 24724 15484
rect 23996 14018 24052 14028
rect 24220 14196 24276 14206
rect 24220 13076 24276 14140
rect 24220 13010 24276 13020
rect 24332 11620 24388 11630
rect 24108 11396 24164 11406
rect 24108 9156 24164 11340
rect 24332 9380 24388 11564
rect 24556 11396 24612 11406
rect 24556 11172 24612 11340
rect 24556 11106 24612 11116
rect 25004 10052 25060 20412
rect 26012 19236 26068 21644
rect 25116 16436 25172 16446
rect 25116 13188 25172 16380
rect 26012 15428 26068 19180
rect 26012 15362 26068 15372
rect 25116 13122 25172 13132
rect 25004 9986 25060 9996
rect 25340 10836 25396 10846
rect 24332 9314 24388 9324
rect 24108 6804 24164 9100
rect 25340 7588 25396 10780
rect 25788 10724 25844 10734
rect 25788 7700 25844 10668
rect 26348 10612 26404 10622
rect 25788 7634 25844 7644
rect 26124 9268 26180 9278
rect 24108 6738 24164 6748
rect 24444 6804 24500 6814
rect 24444 4452 24500 6748
rect 25340 5572 25396 7532
rect 26124 7140 26180 9212
rect 26124 7074 26180 7084
rect 26348 8036 26404 10556
rect 26572 9268 26628 30828
rect 35168 30604 35488 32116
rect 28700 30548 28756 30558
rect 27580 29540 27636 29550
rect 26684 22372 26740 22382
rect 26684 21140 26740 22316
rect 26684 21074 26740 21084
rect 26684 16324 26740 16334
rect 26684 13524 26740 16268
rect 26684 13458 26740 13468
rect 27356 12180 27412 12190
rect 27356 11844 27412 12124
rect 27580 12180 27636 29484
rect 28700 24836 28756 30492
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 28700 24770 28756 24780
rect 28812 26964 28868 26974
rect 27580 12114 27636 12124
rect 27692 18340 27748 18350
rect 27356 11778 27412 11788
rect 26572 9202 26628 9212
rect 25340 5506 25396 5516
rect 24444 4228 24500 4396
rect 24444 4162 24500 4172
rect 26348 4116 26404 7980
rect 26348 4050 26404 4060
rect 27692 1540 27748 18284
rect 28140 14980 28196 14990
rect 28140 12516 28196 14924
rect 28140 12450 28196 12460
rect 28140 5348 28196 5358
rect 28140 5124 28196 5292
rect 28140 5058 28196 5068
rect 28812 3668 28868 26908
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 31836 25284 31892 25294
rect 31612 23828 31668 23838
rect 31612 23604 31668 23772
rect 31612 23538 31668 23548
rect 31500 15652 31556 15662
rect 31500 12628 31556 15596
rect 31500 12562 31556 12572
rect 31836 10724 31892 25228
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 31948 20692 32004 20702
rect 31948 20468 32004 20636
rect 31948 20402 32004 20412
rect 31836 10658 31892 10668
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 28812 3602 28868 3612
rect 29148 10500 29204 10510
rect 29148 2772 29204 10444
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 36988 11844 37044 11854
rect 36988 10052 37044 11788
rect 36988 9986 37044 9996
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 43708 8372 43764 8382
rect 43708 8148 43764 8316
rect 43708 8082 43764 8092
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
rect 29148 2706 29204 2716
rect 27692 1474 27748 1484
rect 23884 1362 23940 1372
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1442_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6160 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1443_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1444_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6832 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1445_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1446_
timestamp 1698431365
transform 1 0 13776 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1447_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14784 0 1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1448_
timestamp 1698431365
transform 1 0 4592 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1449_
timestamp 1698431365
transform -1 0 5376 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1450_
timestamp 1698431365
transform -1 0 5264 0 1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1451_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6384 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1452_
timestamp 1698431365
transform 1 0 7280 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1453_
timestamp 1698431365
transform 1 0 8288 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1454_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 12992 0 1 17248
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1455_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16800 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1456_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25984 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1457_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1458_
timestamp 1698431365
transform -1 0 8624 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1459_
timestamp 1698431365
transform 1 0 7952 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1460_
timestamp 1698431365
transform 1 0 6832 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1461_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9072 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1462_
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1463_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10304 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1464_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 14672 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1465_
timestamp 1698431365
transform -1 0 12320 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1466_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6720 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1467_
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1468_
timestamp 1698431365
transform -1 0 25984 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1469_
timestamp 1698431365
transform 1 0 30016 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1470_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1471_
timestamp 1698431365
transform 1 0 7952 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1472_
timestamp 1698431365
transform -1 0 11424 0 -1 25088
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1473_
timestamp 1698431365
transform 1 0 16240 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1474_
timestamp 1698431365
transform 1 0 24416 0 1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1475_
timestamp 1698431365
transform 1 0 27440 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1476_
timestamp 1698431365
transform 1 0 27888 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1477_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25760 0 1 25088
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1478_
timestamp 1698431365
transform 1 0 29008 0 -1 26656
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1479_
timestamp 1698431365
transform 1 0 31472 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1480_
timestamp 1698431365
transform 1 0 35952 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1481_
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1482_
timestamp 1698431365
transform 1 0 38080 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1483_
timestamp 1698431365
transform -1 0 9184 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1484_
timestamp 1698431365
transform 1 0 6496 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1485_
timestamp 1698431365
transform 1 0 7168 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1486_
timestamp 1698431365
transform 1 0 8288 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1487_
timestamp 1698431365
transform 1 0 11872 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1488_
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1489_
timestamp 1698431365
transform -1 0 13328 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1490_
timestamp 1698431365
transform -1 0 7280 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1491_
timestamp 1698431365
transform 1 0 7056 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1492_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10416 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1493_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12208 0 -1 50176
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1494_
timestamp 1698431365
transform 1 0 21168 0 1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1495_
timestamp 1698431365
transform 1 0 6720 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1496_
timestamp 1698431365
transform 1 0 14560 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1497_
timestamp 1698431365
transform -1 0 9184 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1498_
timestamp 1698431365
transform 1 0 8064 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1499_
timestamp 1698431365
transform 1 0 9072 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1500_
timestamp 1698431365
transform 1 0 8176 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1501_
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1502_
timestamp 1698431365
transform 1 0 6496 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1503_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9744 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1504_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 24080 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1505_
timestamp 1698431365
transform -1 0 23296 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1506_
timestamp 1698431365
transform 1 0 13440 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1507_
timestamp 1698431365
transform -1 0 14896 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1508_
timestamp 1698431365
transform 1 0 24416 0 -1 56448
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1509_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 25984 0 1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1510_
timestamp 1698431365
transform -1 0 23744 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1511_
timestamp 1698431365
transform 1 0 13888 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1512_
timestamp 1698431365
transform 1 0 21168 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1513_
timestamp 1698431365
transform 1 0 14896 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1514_
timestamp 1698431365
transform 1 0 15792 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1515_
timestamp 1698431365
transform 1 0 9408 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1516_
timestamp 1698431365
transform 1 0 5824 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1517_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8400 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1518_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18592 0 -1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1519_
timestamp 1698431365
transform -1 0 31808 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1520_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30016 0 -1 47040
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1521_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 37968 0 -1 37632
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1522_
timestamp 1698431365
transform 1 0 38976 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1523_
timestamp 1698431365
transform 1 0 32256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1524_
timestamp 1698431365
transform -1 0 35056 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1525_
timestamp 1698431365
transform 1 0 36400 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1526_
timestamp 1698431365
transform -1 0 35504 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1527_
timestamp 1698431365
transform 1 0 41216 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1528_
timestamp 1698431365
transform 1 0 36624 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1529_
timestamp 1698431365
transform 1 0 37184 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1530_
timestamp 1698431365
transform -1 0 38864 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1531_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36960 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1532_
timestamp 1698431365
transform -1 0 35840 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1533_
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1534_
timestamp 1698431365
transform 1 0 38640 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1535_
timestamp 1698431365
transform -1 0 39536 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1536_
timestamp 1698431365
transform 1 0 39424 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1537_
timestamp 1698431365
transform 1 0 37968 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1538_
timestamp 1698431365
transform -1 0 42224 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1539_
timestamp 1698431365
transform 1 0 38416 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1540_
timestamp 1698431365
transform 1 0 39312 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1541_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1542_
timestamp 1698431365
transform 1 0 38192 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1543_
timestamp 1698431365
transform -1 0 39984 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1544_
timestamp 1698431365
transform -1 0 39088 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1545_
timestamp 1698431365
transform -1 0 34608 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1546_
timestamp 1698431365
transform 1 0 8064 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1547_
timestamp 1698431365
transform 1 0 8848 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1548_
timestamp 1698431365
transform 1 0 7168 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1549_
timestamp 1698431365
transform 1 0 7728 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1550_
timestamp 1698431365
transform 1 0 9296 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1551_
timestamp 1698431365
transform 1 0 15568 0 1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1552_
timestamp 1698431365
transform 1 0 29008 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1553_
timestamp 1698431365
transform -1 0 7504 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1554_
timestamp 1698431365
transform 1 0 7504 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1555_
timestamp 1698431365
transform 1 0 10640 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1556_
timestamp 1698431365
transform -1 0 11424 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1557_
timestamp 1698431365
transform 1 0 10192 0 1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1558_
timestamp 1698431365
transform 1 0 24192 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1559_
timestamp 1698431365
transform -1 0 29904 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1560_
timestamp 1698431365
transform 1 0 20048 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1561_
timestamp 1698431365
transform 1 0 10080 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1562_
timestamp 1698431365
transform 1 0 15456 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1563_
timestamp 1698431365
transform 1 0 13328 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1564_
timestamp 1698431365
transform 1 0 7728 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1565_
timestamp 1698431365
transform 1 0 11536 0 1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1566_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16016 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1567_
timestamp 1698431365
transform 1 0 30128 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1568_
timestamp 1698431365
transform 1 0 17696 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1569_
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1570_
timestamp 1698431365
transform 1 0 18592 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1571_
timestamp 1698431365
transform 1 0 20944 0 -1 48608
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1572_
timestamp 1698431365
transform 1 0 7504 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1573_
timestamp 1698431365
transform 1 0 14896 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1574_
timestamp 1698431365
transform 1 0 24080 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1575_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31136 0 -1 50176
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1576_
timestamp 1698431365
transform 1 0 25424 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1577_
timestamp 1698431365
transform 1 0 31808 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1578_
timestamp 1698431365
transform -1 0 33488 0 1 53312
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1579_
timestamp 1698431365
transform 1 0 9968 0 1 51744
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1580_
timestamp 1698431365
transform 1 0 9744 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1581_
timestamp 1698431365
transform 1 0 25312 0 -1 50176
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1582_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1583_
timestamp 1698431365
transform 1 0 10640 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1584_
timestamp 1698431365
transform 1 0 19376 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1585_
timestamp 1698431365
transform 1 0 12432 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1586_
timestamp 1698431365
transform 1 0 23632 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1587_
timestamp 1698431365
transform -1 0 28336 0 1 43904
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1588_
timestamp 1698431365
transform -1 0 26544 0 -1 54880
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1589_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33712 0 1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1590_
timestamp 1698431365
transform 1 0 46368 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1591_
timestamp 1698431365
transform -1 0 46704 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1592_
timestamp 1698431365
transform 1 0 45584 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1593_
timestamp 1698431365
transform 1 0 48272 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1594_
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1595_
timestamp 1698431365
transform 1 0 18480 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1596_
timestamp 1698431365
transform 1 0 10976 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1597_
timestamp 1698431365
transform 1 0 11984 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1598_
timestamp 1698431365
transform 1 0 6384 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1599_
timestamp 1698431365
transform 1 0 6832 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1600_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7840 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1601_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 13104 0 1 48608
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1602_
timestamp 1698431365
transform 1 0 13328 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1603_
timestamp 1698431365
transform 1 0 14560 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  _1604_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15008 0 -1 37632
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _1605_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _1606_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30240 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1607_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19712 0 1 53312
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1608_
timestamp 1698431365
transform 1 0 7392 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1609_
timestamp 1698431365
transform 1 0 11648 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1610_
timestamp 1698431365
transform -1 0 17360 0 1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1611_
timestamp 1698431365
transform 1 0 17584 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1612_
timestamp 1698431365
transform -1 0 10192 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1613_
timestamp 1698431365
transform 1 0 7056 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1614_
timestamp 1698431365
transform 1 0 8848 0 1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1615_
timestamp 1698431365
transform -1 0 11648 0 -1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1616_
timestamp 1698431365
transform 1 0 18592 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1617_
timestamp 1698431365
transform 1 0 17696 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1618_
timestamp 1698431365
transform -1 0 12768 0 1 51744
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1619_
timestamp 1698431365
transform -1 0 13104 0 1 53312
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1620_
timestamp 1698431365
transform 1 0 17248 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _1621_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17584 0 -1 54880
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1622_
timestamp 1698431365
transform 1 0 47600 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1623_
timestamp 1698431365
transform -1 0 47600 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1624_
timestamp 1698431365
transform 1 0 23632 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1625_
timestamp 1698431365
transform 1 0 16800 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1626_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23296 0 1 54880
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1627_
timestamp 1698431365
transform 1 0 21504 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1628_
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1629_
timestamp 1698431365
transform 1 0 16128 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1630_
timestamp 1698431365
transform 1 0 12544 0 -1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1631_
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1632_
timestamp 1698431365
transform -1 0 14560 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1633_
timestamp 1698431365
transform 1 0 20496 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1634_
timestamp 1698431365
transform 1 0 15568 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1635_
timestamp 1698431365
transform 1 0 19712 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1636_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22736 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1637_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9184 0 1 36064
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1638_
timestamp 1698431365
transform -1 0 10080 0 1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1639_
timestamp 1698431365
transform -1 0 13104 0 1 40768
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1640_
timestamp 1698431365
transform 1 0 14784 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1641_
timestamp 1698431365
transform 1 0 10192 0 -1 53312
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1642_
timestamp 1698431365
transform 1 0 20496 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1643_
timestamp 1698431365
transform -1 0 20944 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1644_
timestamp 1698431365
transform 1 0 19488 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1645_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 50176
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1646_
timestamp 1698431365
transform 1 0 39312 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1647_
timestamp 1698431365
transform 1 0 40544 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1648_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 39200 0 1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1649_
timestamp 1698431365
transform 1 0 41216 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1650_
timestamp 1698431365
transform 1 0 39872 0 1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1651_
timestamp 1698431365
transform 1 0 41216 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1652_
timestamp 1698431365
transform 1 0 47264 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1653_
timestamp 1698431365
transform 1 0 48608 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1654_
timestamp 1698431365
transform -1 0 30912 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1655_
timestamp 1698431365
transform -1 0 32928 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  _1656_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29456 0 1 54880
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1657_
timestamp 1698431365
transform 1 0 18592 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1658_
timestamp 1698431365
transform 1 0 19600 0 -1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1659_
timestamp 1698431365
transform -1 0 28896 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1660_
timestamp 1698431365
transform 1 0 26992 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1661_
timestamp 1698431365
transform 1 0 14448 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1662_
timestamp 1698431365
transform 1 0 15344 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1663_
timestamp 1698431365
transform -1 0 27104 0 -1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1664_
timestamp 1698431365
transform 1 0 10752 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1665_
timestamp 1698431365
transform 1 0 25872 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1666_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31136 0 -1 50176
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1667_
timestamp 1698431365
transform 1 0 18928 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1668_
timestamp 1698431365
transform 1 0 16352 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1669_
timestamp 1698431365
transform 1 0 19152 0 -1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1670_
timestamp 1698431365
transform 1 0 16688 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1671_
timestamp 1698431365
transform -1 0 24864 0 -1 54880
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_4  _1672_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26880 0 -1 54880
box -86 -86 5798 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1673_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 43344 0 -1 54880
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1674_
timestamp 1698431365
transform 1 0 38416 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1675_
timestamp 1698431365
transform -1 0 38416 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1676_
timestamp 1698431365
transform 1 0 23968 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1677_
timestamp 1698431365
transform 1 0 20048 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1678_
timestamp 1698431365
transform -1 0 18928 0 -1 51744
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1679_
timestamp 1698431365
transform 1 0 22064 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1680_
timestamp 1698431365
transform 1 0 21168 0 1 53312
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1681_
timestamp 1698431365
transform 1 0 7168 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1682_
timestamp 1698431365
transform 1 0 9520 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1683_
timestamp 1698431365
transform 1 0 19712 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1684_
timestamp 1698431365
transform 1 0 7168 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1685_
timestamp 1698431365
transform 1 0 15008 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1686_
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1687_
timestamp 1698431365
transform 1 0 16128 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1688_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1689_
timestamp 1698431365
transform 1 0 22736 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1690_
timestamp 1698431365
transform 1 0 23184 0 1 48608
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1691_
timestamp 1698431365
transform 1 0 35168 0 1 54880
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1692_
timestamp 1698431365
transform -1 0 20944 0 1 54880
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1693_
timestamp 1698431365
transform 1 0 26880 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1694_
timestamp 1698431365
transform 1 0 13888 0 -1 53312
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1695_
timestamp 1698431365
transform 1 0 22960 0 1 53312
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1696_
timestamp 1698431365
transform 1 0 18256 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1697_
timestamp 1698431365
transform 1 0 18256 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1698_
timestamp 1698431365
transform 1 0 23968 0 1 51744
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__or3_2  _1699_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7840 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1700_
timestamp 1698431365
transform 1 0 10976 0 -1 51744
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1701_
timestamp 1698431365
transform 1 0 13328 0 1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1702_
timestamp 1698431365
transform -1 0 15904 0 -1 51744
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1703_
timestamp 1698431365
transform 1 0 11536 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1704_
timestamp 1698431365
transform -1 0 15456 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1705_
timestamp 1698431365
transform -1 0 17920 0 1 51744
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1706_
timestamp 1698431365
transform -1 0 23072 0 -1 53312
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1707_
timestamp 1698431365
transform -1 0 28672 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1708_
timestamp 1698431365
transform -1 0 39984 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1709_
timestamp 1698431365
transform 1 0 37856 0 -1 54880
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1710_
timestamp 1698431365
transform -1 0 46928 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1711_
timestamp 1698431365
transform 1 0 44016 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1712_
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _1713_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7168 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1714_
timestamp 1698431365
transform 1 0 13664 0 1 42336
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1715_
timestamp 1698431365
transform 1 0 16352 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1716_
timestamp 1698431365
transform -1 0 19152 0 1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1717_
timestamp 1698431365
transform 1 0 10080 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1718_
timestamp 1698431365
transform -1 0 20496 0 -1 51744
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1719_
timestamp 1698431365
transform -1 0 20496 0 1 39200
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1720_
timestamp 1698431365
transform 1 0 20384 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1721_
timestamp 1698431365
transform 1 0 31248 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1722_
timestamp 1698431365
transform 1 0 29680 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1723_
timestamp 1698431365
transform 1 0 32928 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1724_
timestamp 1698431365
transform 1 0 30464 0 1 51744
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1725_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 39536 0 -1 51744
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1726_
timestamp 1698431365
transform -1 0 44016 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1727_
timestamp 1698431365
transform -1 0 38752 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1728_
timestamp 1698431365
transform -1 0 18592 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1729_
timestamp 1698431365
transform 1 0 20048 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1730_
timestamp 1698431365
transform 1 0 23296 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1731_
timestamp 1698431365
transform -1 0 20048 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1732_
timestamp 1698431365
transform 1 0 9072 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1733_
timestamp 1698431365
transform -1 0 15792 0 1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1734_
timestamp 1698431365
transform 1 0 21616 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1735_
timestamp 1698431365
transform 1 0 17920 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1736_
timestamp 1698431365
transform 1 0 21728 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1737_
timestamp 1698431365
transform 1 0 22848 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1738_
timestamp 1698431365
transform 1 0 16128 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1739_
timestamp 1698431365
transform 1 0 24192 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1740_
timestamp 1698431365
transform 1 0 14672 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1741_
timestamp 1698431365
transform 1 0 26544 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1742_
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1743_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28336 0 -1 45472
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1744_
timestamp 1698431365
transform 1 0 33264 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1745_
timestamp 1698431365
transform 1 0 33600 0 1 43904
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1746_
timestamp 1698431365
transform -1 0 32480 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1747_
timestamp 1698431365
transform -1 0 22736 0 1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1748_
timestamp 1698431365
transform 1 0 10416 0 -1 40768
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1749_
timestamp 1698431365
transform -1 0 31248 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1750_
timestamp 1698431365
transform 1 0 35616 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1751_
timestamp 1698431365
transform 1 0 29680 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1752_
timestamp 1698431365
transform 1 0 30576 0 -1 51744
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1753_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 38304 0 1 50176
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1754_
timestamp 1698431365
transform 1 0 40768 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1755_
timestamp 1698431365
transform 1 0 42112 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1756_
timestamp 1698431365
transform 1 0 43008 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1757_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 43344 0 -1 54880
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1758_
timestamp 1698431365
transform 1 0 42896 0 1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1759_
timestamp 1698431365
transform 1 0 44800 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1760_
timestamp 1698431365
transform -1 0 42896 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1761_
timestamp 1698431365
transform 1 0 32928 0 -1 54880
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1762_
timestamp 1698431365
transform 1 0 35056 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1763_
timestamp 1698431365
transform 1 0 37072 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1764_
timestamp 1698431365
transform 1 0 20272 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1765_
timestamp 1698431365
transform -1 0 28784 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1766_
timestamp 1698431365
transform 1 0 21392 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1767_
timestamp 1698431365
transform -1 0 25872 0 -1 51744
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1768_
timestamp 1698431365
transform 1 0 32256 0 1 50176
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1769_
timestamp 1698431365
transform 1 0 23744 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1770_
timestamp 1698431365
transform -1 0 10192 0 1 48608
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1771_
timestamp 1698431365
transform 1 0 12208 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _1772_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23632 0 1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1773_
timestamp 1698431365
transform -1 0 14672 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1774_
timestamp 1698431365
transform 1 0 15120 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1775_
timestamp 1698431365
transform 1 0 19712 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1776_
timestamp 1698431365
transform 1 0 21168 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1777_
timestamp 1698431365
transform 1 0 14448 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1778_
timestamp 1698431365
transform 1 0 23744 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1779_
timestamp 1698431365
transform 1 0 24080 0 -1 45472
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1780_
timestamp 1698431365
transform 1 0 25088 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1781_
timestamp 1698431365
transform 1 0 34160 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1782_
timestamp 1698431365
transform 1 0 35056 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1783_
timestamp 1698431365
transform 1 0 35840 0 -1 54880
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1784_
timestamp 1698431365
transform 1 0 47488 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1785_
timestamp 1698431365
transform -1 0 42224 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1786_
timestamp 1698431365
transform 1 0 27440 0 -1 53312
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1787_
timestamp 1698431365
transform 1 0 40768 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1788_
timestamp 1698431365
transform 1 0 7728 0 -1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1789_
timestamp 1698431365
transform 1 0 11984 0 -1 43904
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1790_
timestamp 1698431365
transform -1 0 17024 0 -1 48608
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1791_
timestamp 1698431365
transform 1 0 12208 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1792_
timestamp 1698431365
transform 1 0 12768 0 -1 42336
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1793_
timestamp 1698431365
transform -1 0 12208 0 -1 48608
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1794_
timestamp 1698431365
transform -1 0 15008 0 1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1795_
timestamp 1698431365
transform 1 0 13328 0 1 47040
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1796_
timestamp 1698431365
transform 1 0 18144 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1797_
timestamp 1698431365
transform 1 0 30352 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1798_
timestamp 1698431365
transform -1 0 20720 0 1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1799_
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1800_
timestamp 1698431365
transform 1 0 37184 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1801_
timestamp 1698431365
transform 1 0 38192 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1802_
timestamp 1698431365
transform 1 0 39648 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1803_
timestamp 1698431365
transform -1 0 40432 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1804_
timestamp 1698431365
transform 1 0 40544 0 1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1805_
timestamp 1698431365
transform 1 0 39312 0 1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1806_
timestamp 1698431365
transform 1 0 42560 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1807_
timestamp 1698431365
transform 1 0 43344 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1808_
timestamp 1698431365
transform -1 0 20944 0 1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1809_
timestamp 1698431365
transform 1 0 20048 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1810_
timestamp 1698431365
transform -1 0 28672 0 1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1811_
timestamp 1698431365
transform -1 0 23744 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1812_
timestamp 1698431365
transform 1 0 14672 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1813_
timestamp 1698431365
transform 1 0 22400 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1814_
timestamp 1698431365
transform 1 0 9856 0 -1 45472
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1815_
timestamp 1698431365
transform -1 0 18704 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1816_
timestamp 1698431365
transform 1 0 21168 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1817_
timestamp 1698431365
transform 1 0 14336 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1818_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1819_
timestamp 1698431365
transform 1 0 22064 0 -1 47040
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1820_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26768 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1821_
timestamp 1698431365
transform 1 0 42336 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1822_
timestamp 1698431365
transform 1 0 43120 0 1 51744
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1823_
timestamp 1698431365
transform -1 0 45584 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1824_
timestamp 1698431365
transform 1 0 45248 0 -1 53312
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1825_
timestamp 1698431365
transform 1 0 49728 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_2  _1826_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 47712 0 1 54880
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1827_
timestamp 1698431365
transform 1 0 50960 0 1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1828_
timestamp 1698431365
transform 1 0 52528 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1829_
timestamp 1698431365
transform 1 0 45584 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1830_
timestamp 1698431365
transform 1 0 47152 0 1 53312
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1831_
timestamp 1698431365
transform 1 0 36848 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1832_
timestamp 1698431365
transform 1 0 35952 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1833_
timestamp 1698431365
transform 1 0 6944 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1834_
timestamp 1698431365
transform 1 0 15904 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1835_
timestamp 1698431365
transform 1 0 28224 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1836_
timestamp 1698431365
transform -1 0 25872 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1837_
timestamp 1698431365
transform 1 0 28224 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1838_
timestamp 1698431365
transform 1 0 27104 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1839_
timestamp 1698431365
transform -1 0 28224 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1840_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27104 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1841_
timestamp 1698431365
transform -1 0 30016 0 1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1842_
timestamp 1698431365
transform -1 0 26656 0 -1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1843_
timestamp 1698431365
transform 1 0 31360 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1844_
timestamp 1698431365
transform 1 0 32256 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1845_
timestamp 1698431365
transform 1 0 33376 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1846_
timestamp 1698431365
transform 1 0 34272 0 -1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1847_
timestamp 1698431365
transform 1 0 36848 0 1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1848_
timestamp 1698431365
transform 1 0 45472 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1849_
timestamp 1698431365
transform 1 0 10752 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1850_
timestamp 1698431365
transform 1 0 9856 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1851_
timestamp 1698431365
transform -1 0 10416 0 -1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1852_
timestamp 1698431365
transform -1 0 12208 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1853_
timestamp 1698431365
transform 1 0 10304 0 -1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1854_
timestamp 1698431365
transform -1 0 19152 0 -1 50176
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1855_
timestamp 1698431365
transform 1 0 13664 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1856_
timestamp 1698431365
transform -1 0 16016 0 1 40768
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1857_
timestamp 1698431365
transform 1 0 14112 0 -1 47040
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1858_
timestamp 1698431365
transform -1 0 9744 0 1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1859_
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1860_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15904 0 1 43904
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1861_
timestamp 1698431365
transform -1 0 17136 0 1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1862_
timestamp 1698431365
transform 1 0 17136 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1863_
timestamp 1698431365
transform 1 0 43456 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1864_
timestamp 1698431365
transform 1 0 43008 0 1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1865_
timestamp 1698431365
transform 1 0 38976 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1866_
timestamp 1698431365
transform 1 0 19376 0 -1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1867_
timestamp 1698431365
transform 1 0 22176 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1868_
timestamp 1698431365
transform 1 0 21504 0 1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1869_
timestamp 1698431365
transform -1 0 17696 0 1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1870_
timestamp 1698431365
transform 1 0 16128 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1871_
timestamp 1698431365
transform 1 0 18816 0 1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1872_
timestamp 1698431365
transform -1 0 19488 0 1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1873_
timestamp 1698431365
transform 1 0 17248 0 -1 48608
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1874_
timestamp 1698431365
transform 1 0 38080 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1875_
timestamp 1698431365
transform -1 0 40096 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1876_
timestamp 1698431365
transform 1 0 38976 0 -1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1877_
timestamp 1698431365
transform -1 0 47264 0 -1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1878_
timestamp 1698431365
transform 1 0 46368 0 1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _1879_
timestamp 1698431365
transform 1 0 48272 0 1 50176
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1880_
timestamp 1698431365
transform 1 0 48608 0 -1 51744
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1881_
timestamp 1698431365
transform 1 0 50848 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1882_
timestamp 1698431365
transform 1 0 47264 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1883_
timestamp 1698431365
transform 1 0 47264 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1884_
timestamp 1698431365
transform -1 0 47264 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1885_
timestamp 1698431365
transform 1 0 48608 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1886_
timestamp 1698431365
transform -1 0 51296 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1887_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 51072 0 -1 53312
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1888_
timestamp 1698431365
transform 1 0 53424 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1889_
timestamp 1698431365
transform 1 0 49952 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1890_
timestamp 1698431365
transform 1 0 50512 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1891_
timestamp 1698431365
transform 1 0 27664 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1892_
timestamp 1698431365
transform 1 0 26544 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1893_
timestamp 1698431365
transform 1 0 21616 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1894_
timestamp 1698431365
transform 1 0 26768 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1895_
timestamp 1698431365
transform 1 0 24304 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1896_
timestamp 1698431365
transform 1 0 25200 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1897_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26208 0 -1 42336
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1898_
timestamp 1698431365
transform 1 0 29344 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1899_
timestamp 1698431365
transform 1 0 27216 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1900_
timestamp 1698431365
transform 1 0 29008 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1901_
timestamp 1698431365
transform -1 0 29344 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1902_
timestamp 1698431365
transform -1 0 29568 0 -1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1903_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1904_
timestamp 1698431365
transform 1 0 30240 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1905_
timestamp 1698431365
transform 1 0 33376 0 -1 51744
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1906_
timestamp 1698431365
transform -1 0 39200 0 -1 51744
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1907_
timestamp 1698431365
transform 1 0 38080 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1908_
timestamp 1698431365
transform 1 0 37408 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1909_
timestamp 1698431365
transform -1 0 46368 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1910_
timestamp 1698431365
transform -1 0 46256 0 1 48608
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1911_
timestamp 1698431365
transform 1 0 19488 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1912_
timestamp 1698431365
transform -1 0 17920 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1913_
timestamp 1698431365
transform 1 0 13104 0 -1 40768
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1914_
timestamp 1698431365
transform -1 0 13552 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _1915_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 45472
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1916_
timestamp 1698431365
transform 1 0 15904 0 1 45472
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1917_
timestamp 1698431365
transform -1 0 24192 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1918_
timestamp 1698431365
transform 1 0 44688 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1919_
timestamp 1698431365
transform 1 0 45024 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1920_
timestamp 1698431365
transform -1 0 46480 0 -1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1921_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37520 0 -1 48608
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1922_
timestamp 1698431365
transform 1 0 40096 0 1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1923_
timestamp 1698431365
transform 1 0 22512 0 -1 42336
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1924_
timestamp 1698431365
transform -1 0 22288 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1925_
timestamp 1698431365
transform 1 0 22176 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1926_
timestamp 1698431365
transform -1 0 11648 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1927_
timestamp 1698431365
transform -1 0 23632 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1928_
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1929_
timestamp 1698431365
transform -1 0 21728 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1930_
timestamp 1698431365
transform -1 0 22512 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1931_
timestamp 1698431365
transform 1 0 27888 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1932_
timestamp 1698431365
transform 1 0 38416 0 1 43904
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1933_
timestamp 1698431365
transform 1 0 42224 0 -1 47040
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1934_
timestamp 1698431365
transform 1 0 48608 0 -1 47040
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1935_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 46592 0 1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1936_
timestamp 1698431365
transform 1 0 48832 0 -1 48608
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1937_
timestamp 1698431365
transform 1 0 49616 0 -1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _1938_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 50176 0 -1 50176
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1939_
timestamp 1698431365
transform -1 0 52304 0 1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1940_
timestamp 1698431365
transform 1 0 49952 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1941_
timestamp 1698431365
transform 1 0 51296 0 -1 54880
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1942_
timestamp 1698431365
transform 1 0 52528 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1943_
timestamp 1698431365
transform 1 0 53424 0 1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1944_
timestamp 1698431365
transform 1 0 54544 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1945_
timestamp 1698431365
transform -1 0 52080 0 1 47040
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1946_
timestamp 1698431365
transform 1 0 49840 0 -1 47040
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1947_
timestamp 1698431365
transform 1 0 52864 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1948_
timestamp 1698431365
transform 1 0 24976 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1949_
timestamp 1698431365
transform 1 0 26432 0 1 45472
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1950_
timestamp 1698431365
transform 1 0 29456 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1951_
timestamp 1698431365
transform -1 0 30240 0 1 43904
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1952_
timestamp 1698431365
transform -1 0 27216 0 1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1953_
timestamp 1698431365
transform 1 0 30576 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1954_
timestamp 1698431365
transform -1 0 35616 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1955_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31472 0 1 43904
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1956_
timestamp 1698431365
transform 1 0 35952 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1957_
timestamp 1698431365
transform -1 0 38080 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1958_
timestamp 1698431365
transform 1 0 37072 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1959_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 45472 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1960_
timestamp 1698431365
transform -1 0 20608 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1961_
timestamp 1698431365
transform 1 0 20048 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1962_
timestamp 1698431365
transform 1 0 21168 0 1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1963_
timestamp 1698431365
transform 1 0 19264 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1964_
timestamp 1698431365
transform -1 0 30464 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1965_
timestamp 1698431365
transform 1 0 35504 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1966_
timestamp 1698431365
transform -1 0 36736 0 -1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1967_
timestamp 1698431365
transform 1 0 44800 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1968_
timestamp 1698431365
transform -1 0 45696 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1969_
timestamp 1698431365
transform 1 0 40768 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1970_
timestamp 1698431365
transform 1 0 37296 0 1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1971_
timestamp 1698431365
transform 1 0 30240 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1972_
timestamp 1698431365
transform -1 0 29904 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1973_
timestamp 1698431365
transform -1 0 32368 0 1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1974_
timestamp 1698431365
transform -1 0 19600 0 1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1975_
timestamp 1698431365
transform -1 0 27328 0 1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _1976_
timestamp 1698431365
transform 1 0 23072 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1977_
timestamp 1698431365
transform -1 0 34832 0 -1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1978_
timestamp 1698431365
transform 1 0 33264 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1979_
timestamp 1698431365
transform 1 0 34832 0 -1 48608
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1980_
timestamp 1698431365
transform 1 0 35840 0 -1 47040
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1981_
timestamp 1698431365
transform 1 0 38528 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1982_
timestamp 1698431365
transform 1 0 39648 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1983_
timestamp 1698431365
transform 1 0 34832 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1984_
timestamp 1698431365
transform -1 0 36400 0 1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1985_
timestamp 1698431365
transform -1 0 40544 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1986_
timestamp 1698431365
transform 1 0 39872 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1987_
timestamp 1698431365
transform 1 0 40656 0 1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1988_
timestamp 1698431365
transform 1 0 46480 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1989_
timestamp 1698431365
transform -1 0 47712 0 1 43904
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1990_
timestamp 1698431365
transform -1 0 50064 0 -1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1991_
timestamp 1698431365
transform 1 0 50176 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1992_
timestamp 1698431365
transform 1 0 52528 0 1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1993_
timestamp 1698431365
transform 1 0 51520 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1994_
timestamp 1698431365
transform -1 0 53424 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1995_
timestamp 1698431365
transform 1 0 53424 0 1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1996_
timestamp 1698431365
transform 1 0 54768 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1997_
timestamp 1698431365
transform 1 0 50064 0 -1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1998_
timestamp 1698431365
transform 1 0 36288 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _1999_
timestamp 1698431365
transform 1 0 37632 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2000_
timestamp 1698431365
transform -1 0 33600 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2001_
timestamp 1698431365
transform 1 0 22512 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2002_
timestamp 1698431365
transform -1 0 25312 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2003_
timestamp 1698431365
transform 1 0 30464 0 -1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2004_
timestamp 1698431365
transform 1 0 33488 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2005_
timestamp 1698431365
transform -1 0 36176 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2006_
timestamp 1698431365
transform 1 0 34384 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2007_
timestamp 1698431365
transform 1 0 34496 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2008_
timestamp 1698431365
transform 1 0 37632 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2009_
timestamp 1698431365
transform -1 0 46368 0 1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2010_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2011_
timestamp 1698431365
transform 1 0 26208 0 1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2012_
timestamp 1698431365
transform 1 0 27216 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2013_
timestamp 1698431365
transform -1 0 29344 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2014_
timestamp 1698431365
transform -1 0 28560 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2015_
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2016_
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2017_
timestamp 1698431365
transform -1 0 29680 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _2018_
timestamp 1698431365
transform 1 0 26992 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2019_
timestamp 1698431365
transform 1 0 44688 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2020_
timestamp 1698431365
transform 1 0 41216 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2021_
timestamp 1698431365
transform -1 0 34832 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2022_
timestamp 1698431365
transform -1 0 35056 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2023_
timestamp 1698431365
transform -1 0 23184 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2024_
timestamp 1698431365
transform -1 0 23856 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2025_
timestamp 1698431365
transform -1 0 22624 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai33_1  _2026_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22848 0 1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2027_
timestamp 1698431365
transform 1 0 35616 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2028_
timestamp 1698431365
transform -1 0 35616 0 -1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2029_
timestamp 1698431365
transform 1 0 38528 0 1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2030_
timestamp 1698431365
transform 1 0 41216 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2031_
timestamp 1698431365
transform -1 0 42672 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2032_
timestamp 1698431365
transform 1 0 41552 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2033_
timestamp 1698431365
transform 1 0 45472 0 1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2034_
timestamp 1698431365
transform 1 0 44464 0 -1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2035_
timestamp 1698431365
transform -1 0 42224 0 -1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2036_
timestamp 1698431365
transform -1 0 42336 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2037_
timestamp 1698431365
transform -1 0 48048 0 -1 42336
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2038_
timestamp 1698431365
transform 1 0 47824 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2039_
timestamp 1698431365
transform -1 0 49504 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2040_
timestamp 1698431365
transform 1 0 51184 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2041_
timestamp 1698431365
transform 1 0 52528 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2042_
timestamp 1698431365
transform -1 0 56224 0 -1 50176
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2043_
timestamp 1698431365
transform -1 0 52864 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2044_
timestamp 1698431365
transform 1 0 51632 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2045_
timestamp 1698431365
transform -1 0 53984 0 -1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2046_
timestamp 1698431365
transform 1 0 53424 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2047_
timestamp 1698431365
transform 1 0 54096 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2048_
timestamp 1698431365
transform 1 0 55440 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2049_
timestamp 1698431365
transform 1 0 46032 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2050_
timestamp 1698431365
transform 1 0 45920 0 -1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2051_
timestamp 1698431365
transform 1 0 47152 0 1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2052_
timestamp 1698431365
transform -1 0 35392 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2053_
timestamp 1698431365
transform -1 0 33600 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2054_
timestamp 1698431365
transform 1 0 29232 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2055_
timestamp 1698431365
transform -1 0 32592 0 -1 37632
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2056_
timestamp 1698431365
transform -1 0 35616 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2057_
timestamp 1698431365
transform 1 0 34048 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2058_
timestamp 1698431365
transform 1 0 35056 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2059_
timestamp 1698431365
transform 1 0 34720 0 1 37632
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2060_
timestamp 1698431365
transform 1 0 38080 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2061_
timestamp 1698431365
transform 1 0 30464 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2062_
timestamp 1698431365
transform -1 0 32816 0 1 40768
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2063_
timestamp 1698431365
transform 1 0 26096 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2064_
timestamp 1698431365
transform 1 0 26768 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2065_
timestamp 1698431365
transform -1 0 32368 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2066_
timestamp 1698431365
transform -1 0 31808 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2067_
timestamp 1698431365
transform 1 0 25872 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _2068_
timestamp 1698431365
transform 1 0 31360 0 1 37632
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2069_
timestamp 1698431365
transform 1 0 42896 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2070_
timestamp 1698431365
transform -1 0 42896 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2071_
timestamp 1698431365
transform -1 0 45360 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2072_
timestamp 1698431365
transform -1 0 28672 0 1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2073_
timestamp 1698431365
transform -1 0 26768 0 -1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2074_
timestamp 1698431365
transform -1 0 31136 0 -1 39200
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2075_
timestamp 1698431365
transform 1 0 44016 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _2076_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42000 0 1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2077_
timestamp 1698431365
transform -1 0 47936 0 -1 39200
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2078_
timestamp 1698431365
transform -1 0 47152 0 1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2079_
timestamp 1698431365
transform 1 0 44912 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2080_
timestamp 1698431365
transform -1 0 49392 0 1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2081_
timestamp 1698431365
transform 1 0 48608 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2082_
timestamp 1698431365
transform -1 0 49728 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2083_
timestamp 1698431365
transform 1 0 51184 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2084_
timestamp 1698431365
transform -1 0 52080 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2085_
timestamp 1698431365
transform -1 0 53200 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2086_
timestamp 1698431365
transform 1 0 51184 0 -1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2087_
timestamp 1698431365
transform -1 0 54320 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2088_
timestamp 1698431365
transform 1 0 54320 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2089_
timestamp 1698431365
transform -1 0 57120 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2090_
timestamp 1698431365
transform 1 0 53200 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2091_
timestamp 1698431365
transform 1 0 50400 0 -1 40768
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2092_
timestamp 1698431365
transform 1 0 52304 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2093_
timestamp 1698431365
transform 1 0 53200 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2094_
timestamp 1698431365
transform 1 0 51856 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2095_
timestamp 1698431365
transform 1 0 53200 0 1 43904
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2096_
timestamp 1698431365
transform -1 0 51520 0 1 39200
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2097_
timestamp 1698431365
transform 1 0 29120 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2098_
timestamp 1698431365
transform 1 0 29792 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2099_
timestamp 1698431365
transform 1 0 29344 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2100_
timestamp 1698431365
transform 1 0 28336 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2101_
timestamp 1698431365
transform -1 0 32704 0 -1 45472
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _2102_
timestamp 1698431365
transform -1 0 33600 0 1 45472
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2103_
timestamp 1698431365
transform 1 0 41104 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2104_
timestamp 1698431365
transform 1 0 41216 0 -1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2105_
timestamp 1698431365
transform 1 0 42112 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2106_
timestamp 1698431365
transform 1 0 42336 0 -1 43904
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2107_
timestamp 1698431365
transform 1 0 43568 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2108_
timestamp 1698431365
transform 1 0 31360 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2109_
timestamp 1698431365
transform 1 0 32256 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2110_
timestamp 1698431365
transform 1 0 31808 0 1 39200
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2111_
timestamp 1698431365
transform 1 0 32928 0 1 42336
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2112_
timestamp 1698431365
transform -1 0 43792 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2113_
timestamp 1698431365
transform 1 0 44688 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2114_
timestamp 1698431365
transform 1 0 44688 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2115_
timestamp 1698431365
transform -1 0 49616 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2116_
timestamp 1698431365
transform 1 0 49504 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2117_
timestamp 1698431365
transform -1 0 35840 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2118_
timestamp 1698431365
transform -1 0 28448 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2119_
timestamp 1698431365
transform -1 0 25648 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2120_
timestamp 1698431365
transform 1 0 26880 0 -1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2121_
timestamp 1698431365
transform 1 0 37520 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2122_
timestamp 1698431365
transform -1 0 39648 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2123_
timestamp 1698431365
transform 1 0 49616 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2124_
timestamp 1698431365
transform 1 0 50736 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2125_
timestamp 1698431365
transform 1 0 53536 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2126_
timestamp 1698431365
transform -1 0 55552 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2127_
timestamp 1698431365
transform 1 0 54096 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2128_
timestamp 1698431365
transform -1 0 57568 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _2129_
timestamp 1698431365
transform 1 0 49280 0 1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2130_
timestamp 1698431365
transform -1 0 51856 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2131_
timestamp 1698431365
transform -1 0 34384 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2132_
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2133_
timestamp 1698431365
transform 1 0 32592 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2134_
timestamp 1698431365
transform 1 0 34384 0 -1 34496
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2135_
timestamp 1698431365
transform 1 0 37856 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2136_
timestamp 1698431365
transform 1 0 37968 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2137_
timestamp 1698431365
transform 1 0 28560 0 -1 37632
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2138_
timestamp 1698431365
transform 1 0 30576 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2139_
timestamp 1698431365
transform 1 0 31248 0 1 36064
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2140_
timestamp 1698431365
transform -1 0 36288 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2141_
timestamp 1698431365
transform 1 0 41888 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2142_
timestamp 1698431365
transform 1 0 40992 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2143_
timestamp 1698431365
transform -1 0 46928 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2144_
timestamp 1698431365
transform 1 0 42112 0 1 37632
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2145_
timestamp 1698431365
transform 1 0 33824 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2146_
timestamp 1698431365
transform 1 0 35840 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2147_
timestamp 1698431365
transform 1 0 44016 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2148_
timestamp 1698431365
transform 1 0 44576 0 -1 37632
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2149_
timestamp 1698431365
transform 1 0 46928 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2150_
timestamp 1698431365
transform 1 0 48608 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2151_
timestamp 1698431365
transform -1 0 50960 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _2152_
timestamp 1698431365
transform 1 0 50960 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2153_
timestamp 1698431365
transform -1 0 54544 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2154_
timestamp 1698431365
transform -1 0 54432 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2155_
timestamp 1698431365
transform 1 0 54096 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2156_
timestamp 1698431365
transform 1 0 54096 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2157_
timestamp 1698431365
transform 1 0 55552 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2158_
timestamp 1698431365
transform -1 0 32592 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2159_
timestamp 1698431365
transform -1 0 32704 0 -1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2160_
timestamp 1698431365
transform 1 0 33152 0 1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2161_
timestamp 1698431365
transform 1 0 42336 0 1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2162_
timestamp 1698431365
transform 1 0 42000 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2163_
timestamp 1698431365
transform 1 0 43456 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2164_
timestamp 1698431365
transform -1 0 34608 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2165_
timestamp 1698431365
transform 1 0 44688 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2166_
timestamp 1698431365
transform 1 0 44688 0 1 36064
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2167_
timestamp 1698431365
transform 1 0 46816 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2168_
timestamp 1698431365
transform 1 0 47376 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2169_
timestamp 1698431365
transform 1 0 47824 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2170_
timestamp 1698431365
transform -1 0 37744 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2171_
timestamp 1698431365
transform 1 0 36064 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2172_
timestamp 1698431365
transform -1 0 38976 0 1 34496
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2173_
timestamp 1698431365
transform 1 0 44912 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2174_
timestamp 1698431365
transform 1 0 48496 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2175_
timestamp 1698431365
transform 1 0 48048 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2176_
timestamp 1698431365
transform 1 0 51184 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2177_
timestamp 1698431365
transform 1 0 47488 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2178_
timestamp 1698431365
transform 1 0 48384 0 1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _2179_
timestamp 1698431365
transform 1 0 52192 0 -1 34496
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2180_
timestamp 1698431365
transform 1 0 52976 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2181_
timestamp 1698431365
transform -1 0 54096 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2182_
timestamp 1698431365
transform -1 0 54096 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2183_
timestamp 1698431365
transform 1 0 54096 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2184_
timestamp 1698431365
transform 1 0 53872 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2185_
timestamp 1698431365
transform 1 0 55104 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2186_
timestamp 1698431365
transform 1 0 29792 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _2187_
timestamp 1698431365
transform 1 0 29792 0 1 34496
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2188_
timestamp 1698431365
transform 1 0 41104 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2189_
timestamp 1698431365
transform 1 0 41104 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2190_
timestamp 1698431365
transform 1 0 42448 0 -1 36064
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2191_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 44688 0 1 32928
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2192_
timestamp 1698431365
transform -1 0 50288 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2193_
timestamp 1698431365
transform 1 0 49392 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2194_
timestamp 1698431365
transform 1 0 50512 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2195_
timestamp 1698431365
transform -1 0 53648 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2196_
timestamp 1698431365
transform 1 0 52528 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2197_
timestamp 1698431365
transform 1 0 53872 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2198_
timestamp 1698431365
transform 1 0 46704 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2199_
timestamp 1698431365
transform -1 0 46704 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2200_
timestamp 1698431365
transform 1 0 46368 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2201_
timestamp 1698431365
transform 1 0 51744 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2202_
timestamp 1698431365
transform 1 0 52528 0 1 34496
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2203_
timestamp 1698431365
transform 1 0 50512 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2204_
timestamp 1698431365
transform 1 0 48608 0 1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2205_
timestamp 1698431365
transform 1 0 49616 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2206_
timestamp 1698431365
transform -1 0 50064 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _2207_
timestamp 1698431365
transform -1 0 49616 0 1 34496
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2208_
timestamp 1698431365
transform 1 0 44688 0 1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2209_
timestamp 1698431365
transform 1 0 46032 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2210_
timestamp 1698431365
transform -1 0 28784 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2211_
timestamp 1698431365
transform -1 0 27776 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2212_
timestamp 1698431365
transform 1 0 27664 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2213_
timestamp 1698431365
transform -1 0 28784 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2214_
timestamp 1698431365
transform 1 0 8848 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2215_
timestamp 1698431365
transform 1 0 8848 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2216_
timestamp 1698431365
transform 1 0 10192 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2217_
timestamp 1698431365
transform -1 0 12768 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2218_
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2219_
timestamp 1698431365
transform 1 0 7616 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2220_
timestamp 1698431365
transform 1 0 7056 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2221_
timestamp 1698431365
transform 1 0 7952 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _2222_
timestamp 1698431365
transform -1 0 11984 0 -1 26656
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2223_
timestamp 1698431365
transform 1 0 10192 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2224_
timestamp 1698431365
transform 1 0 9968 0 -1 18816
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2225_
timestamp 1698431365
transform 1 0 10640 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2226_
timestamp 1698431365
transform -1 0 8848 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2227_
timestamp 1698431365
transform 1 0 7616 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2228_
timestamp 1698431365
transform 1 0 12544 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2229_
timestamp 1698431365
transform 1 0 5936 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2230_
timestamp 1698431365
transform 1 0 11424 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2231_
timestamp 1698431365
transform -1 0 13104 0 1 23520
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2232_
timestamp 1698431365
transform -1 0 9632 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _2233_
timestamp 1698431365
transform 1 0 10304 0 1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _2234_
timestamp 1698431365
transform 1 0 11536 0 -1 20384
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2235_
timestamp 1698431365
transform 1 0 5936 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2236_
timestamp 1698431365
transform 1 0 7952 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2237_
timestamp 1698431365
transform 1 0 11648 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2238_
timestamp 1698431365
transform 1 0 16016 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2239_
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2240_
timestamp 1698431365
transform 1 0 7952 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2241_
timestamp 1698431365
transform 1 0 4816 0 -1 23520
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2242_
timestamp 1698431365
transform 1 0 17584 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2243_
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2244_
timestamp 1698431365
transform 1 0 18032 0 -1 18816
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2245_
timestamp 1698431365
transform 1 0 27888 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2246_
timestamp 1698431365
transform -1 0 27664 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2247_
timestamp 1698431365
transform -1 0 26880 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2248_
timestamp 1698431365
transform 1 0 24864 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2249_
timestamp 1698431365
transform 1 0 25872 0 1 20384
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2250_
timestamp 1698431365
transform 1 0 42000 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2251_
timestamp 1698431365
transform -1 0 40992 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2252_
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _2253_
timestamp 1698431365
transform 1 0 5264 0 -1 26656
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2254_
timestamp 1698431365
transform -1 0 15792 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2255_
timestamp 1698431365
transform 1 0 13104 0 -1 26656
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2256_
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _2257_
timestamp 1698431365
transform -1 0 27440 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2258_
timestamp 1698431365
transform -1 0 16576 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2259_
timestamp 1698431365
transform -1 0 19152 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2260_
timestamp 1698431365
transform 1 0 18480 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2261_
timestamp 1698431365
transform -1 0 30464 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2262_
timestamp 1698431365
transform 1 0 5712 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2263_
timestamp 1698431365
transform 1 0 5152 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _2264_
timestamp 1698431365
transform 1 0 6384 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2265_
timestamp 1698431365
transform 1 0 7728 0 1 23520
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2266_
timestamp 1698431365
transform 1 0 19376 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _2267_
timestamp 1698431365
transform -1 0 9184 0 -1 20384
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2268_
timestamp 1698431365
transform -1 0 24640 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _2269_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17808 0 -1 23520
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2270_
timestamp 1698431365
transform 1 0 30800 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2271_
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2272_
timestamp 1698431365
transform -1 0 24864 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _2273_
timestamp 1698431365
transform 1 0 10416 0 -1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2274_
timestamp 1698431365
transform 1 0 22960 0 1 26656
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2275_
timestamp 1698431365
transform -1 0 18256 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2276_
timestamp 1698431365
transform 1 0 7056 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2277_
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2278_
timestamp 1698431365
transform -1 0 18144 0 1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2279_
timestamp 1698431365
transform -1 0 7952 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2280_
timestamp 1698431365
transform 1 0 8064 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2281_
timestamp 1698431365
transform -1 0 11088 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2282_
timestamp 1698431365
transform -1 0 12544 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2283_
timestamp 1698431365
transform 1 0 9072 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2284_
timestamp 1698431365
transform 1 0 9520 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2285_
timestamp 1698431365
transform 1 0 7168 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2286_
timestamp 1698431365
transform 1 0 18816 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2287_
timestamp 1698431365
transform 1 0 14448 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2288_
timestamp 1698431365
transform 1 0 16128 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2289_
timestamp 1698431365
transform -1 0 17808 0 1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2290_
timestamp 1698431365
transform -1 0 14560 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2291_
timestamp 1698431365
transform -1 0 13104 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _2292_
timestamp 1698431365
transform -1 0 20608 0 1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _2293_
timestamp 1698431365
transform -1 0 9184 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _2294_
timestamp 1698431365
transform 1 0 18032 0 1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2295_
timestamp 1698431365
transform -1 0 27664 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2296_
timestamp 1698431365
transform 1 0 29904 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2297_
timestamp 1698431365
transform 1 0 25200 0 -1 15680
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2298_
timestamp 1698431365
transform 1 0 16128 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _2299_
timestamp 1698431365
transform 1 0 8512 0 1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2300_
timestamp 1698431365
transform -1 0 18704 0 -1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2301_
timestamp 1698431365
transform -1 0 23408 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2302_
timestamp 1698431365
transform 1 0 11984 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2303_
timestamp 1698431365
transform -1 0 13104 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2304_
timestamp 1698431365
transform 1 0 22960 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2305_
timestamp 1698431365
transform -1 0 29904 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2306_
timestamp 1698431365
transform -1 0 28784 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2307_
timestamp 1698431365
transform 1 0 23968 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _2308_
timestamp 1698431365
transform -1 0 26992 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2309_
timestamp 1698431365
transform 1 0 33936 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2310_
timestamp 1698431365
transform -1 0 42784 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2311_
timestamp 1698431365
transform -1 0 41888 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2312_
timestamp 1698431365
transform 1 0 41888 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2313_
timestamp 1698431365
transform 1 0 45248 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2314_
timestamp 1698431365
transform 1 0 41552 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2315_
timestamp 1698431365
transform -1 0 46144 0 1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2316_
timestamp 1698431365
transform 1 0 45696 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2317_
timestamp 1698431365
transform 1 0 46592 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2318_
timestamp 1698431365
transform 1 0 46256 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2319_
timestamp 1698431365
transform 1 0 47152 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _2320_
timestamp 1698431365
transform 1 0 29680 0 1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2321_
timestamp 1698431365
transform 1 0 8176 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2322_
timestamp 1698431365
transform 1 0 17920 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _2323_
timestamp 1698431365
transform 1 0 10080 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _2324_
timestamp 1698431365
transform 1 0 7168 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _2325_
timestamp 1698431365
transform 1 0 12432 0 -1 23520
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2326_
timestamp 1698431365
transform -1 0 22512 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_2  _2327_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19600 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2328_
timestamp 1698431365
transform 1 0 22288 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2329_
timestamp 1698431365
transform 1 0 17024 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2330_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19600 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2331_
timestamp 1698431365
transform -1 0 26880 0 1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2332_
timestamp 1698431365
transform 1 0 29904 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2333_
timestamp 1698431365
transform -1 0 43680 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2334_
timestamp 1698431365
transform 1 0 43008 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2335_
timestamp 1698431365
transform 1 0 31248 0 1 23520
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _2336_
timestamp 1698431365
transform 1 0 7952 0 1 17248
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _2337_
timestamp 1698431365
transform -1 0 16016 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _2338_
timestamp 1698431365
transform -1 0 7952 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _2339_
timestamp 1698431365
transform 1 0 14112 0 1 23520
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2340_
timestamp 1698431365
transform -1 0 19376 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2341_
timestamp 1698431365
transform -1 0 27888 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2342_
timestamp 1698431365
transform 1 0 25424 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2343_
timestamp 1698431365
transform 1 0 22288 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2344_
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _2345_
timestamp 1698431365
transform -1 0 26768 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2346_
timestamp 1698431365
transform 1 0 31808 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2347_
timestamp 1698431365
transform 1 0 34608 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2348_
timestamp 1698431365
transform -1 0 34160 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2349_
timestamp 1698431365
transform 1 0 23296 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2350_
timestamp 1698431365
transform -1 0 26544 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2351_
timestamp 1698431365
transform -1 0 24864 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2352_
timestamp 1698431365
transform 1 0 6720 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2353_
timestamp 1698431365
transform 1 0 14560 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2354_
timestamp 1698431365
transform -1 0 14784 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2355_
timestamp 1698431365
transform -1 0 9968 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2356_
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2357_
timestamp 1698431365
transform 1 0 15344 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2358_
timestamp 1698431365
transform 1 0 6720 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2359_
timestamp 1698431365
transform 1 0 17248 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2360_
timestamp 1698431365
transform -1 0 22512 0 -1 21952
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2361_
timestamp 1698431365
transform 1 0 16016 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2362_
timestamp 1698431365
transform -1 0 17248 0 1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2363_
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _2364_
timestamp 1698431365
transform 1 0 22736 0 -1 21952
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _2365_
timestamp 1698431365
transform -1 0 7728 0 1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _2366_
timestamp 1698431365
transform 1 0 19152 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2367_
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2368_
timestamp 1698431365
transform -1 0 14896 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2369_
timestamp 1698431365
transform -1 0 23856 0 1 15680
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _2370_
timestamp 1698431365
transform 1 0 10192 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2371_
timestamp 1698431365
transform -1 0 29904 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2372_
timestamp 1698431365
transform 1 0 16016 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2373_
timestamp 1698431365
transform -1 0 26768 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2374_
timestamp 1698431365
transform 1 0 29344 0 1 20384
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2375_
timestamp 1698431365
transform -1 0 20720 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2376_
timestamp 1698431365
transform 1 0 7504 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _2377_
timestamp 1698431365
transform -1 0 7168 0 1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2378_
timestamp 1698431365
transform -1 0 20160 0 1 15680
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2379_
timestamp 1698431365
transform -1 0 22400 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2380_
timestamp 1698431365
transform 1 0 11984 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _2381_
timestamp 1698431365
transform 1 0 13104 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2382_
timestamp 1698431365
transform 1 0 20496 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2383_
timestamp 1698431365
transform -1 0 15232 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2384_
timestamp 1698431365
transform 1 0 17360 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2385_
timestamp 1698431365
transform 1 0 17472 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2386_
timestamp 1698431365
transform 1 0 11424 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2387_
timestamp 1698431365
transform -1 0 16016 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2388_
timestamp 1698431365
transform -1 0 16576 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2389_
timestamp 1698431365
transform -1 0 19824 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2390_
timestamp 1698431365
transform -1 0 28672 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2391_
timestamp 1698431365
transform 1 0 21952 0 1 7840
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2392_
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2393_
timestamp 1698431365
transform -1 0 38416 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2394_
timestamp 1698431365
transform 1 0 35728 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2395_
timestamp 1698431365
transform 1 0 18592 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2396_
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2397_
timestamp 1698431365
transform 1 0 22624 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2398_
timestamp 1698431365
transform 1 0 27216 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2399_
timestamp 1698431365
transform -1 0 31360 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2400_
timestamp 1698431365
transform 1 0 28336 0 -1 20384
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2401_
timestamp 1698431365
transform 1 0 17808 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  _2402_
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2403_
timestamp 1698431365
transform -1 0 11536 0 1 12544
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2404_
timestamp 1698431365
transform 1 0 17696 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2405_
timestamp 1698431365
transform -1 0 22176 0 -1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2406_
timestamp 1698431365
transform -1 0 9072 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2407_
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2408_
timestamp 1698431365
transform -1 0 15456 0 1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2409_
timestamp 1698431365
transform -1 0 23632 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2410_
timestamp 1698431365
transform 1 0 21840 0 1 20384
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2411_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 35504 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2412_
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2413_
timestamp 1698431365
transform 1 0 31360 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2414_
timestamp 1698431365
transform 1 0 34832 0 -1 21952
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2415_
timestamp 1698431365
transform 1 0 34496 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2416_
timestamp 1698431365
transform 1 0 34608 0 1 21952
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2417_
timestamp 1698431365
transform 1 0 44912 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2418_
timestamp 1698431365
transform 1 0 45696 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2419_
timestamp 1698431365
transform 1 0 48832 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2420_
timestamp 1698431365
transform 1 0 44800 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2421_
timestamp 1698431365
transform -1 0 46592 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2422_
timestamp 1698431365
transform -1 0 43344 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2423_
timestamp 1698431365
transform -1 0 43568 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _2424_
timestamp 1698431365
transform 1 0 27888 0 -1 23520
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2425_
timestamp 1698431365
transform 1 0 11872 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2426_
timestamp 1698431365
transform -1 0 20384 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2427_
timestamp 1698431365
transform -1 0 20720 0 1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2428_
timestamp 1698431365
transform 1 0 12096 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2429_
timestamp 1698431365
transform -1 0 18480 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2430_
timestamp 1698431365
transform 1 0 19600 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2431_
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2432_
timestamp 1698431365
transform 1 0 10528 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2433_
timestamp 1698431365
transform 1 0 9632 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _2434_
timestamp 1698431365
transform 1 0 10640 0 -1 17248
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _2435_
timestamp 1698431365
transform -1 0 25760 0 1 25088
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2436_
timestamp 1698431365
transform -1 0 28336 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2437_
timestamp 1698431365
transform 1 0 18816 0 -1 14112
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _2438_
timestamp 1698431365
transform -1 0 22512 0 -1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2439_
timestamp 1698431365
transform 1 0 42560 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2440_
timestamp 1698431365
transform 1 0 45696 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2441_
timestamp 1698431365
transform 1 0 42560 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2442_
timestamp 1698431365
transform -1 0 34608 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2443_
timestamp 1698431365
transform 1 0 34832 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _2444_
timestamp 1698431365
transform 1 0 18032 0 1 23520
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2445_
timestamp 1698431365
transform -1 0 18032 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2446_
timestamp 1698431365
transform 1 0 13776 0 1 25088
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2447_
timestamp 1698431365
transform -1 0 29456 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2448_
timestamp 1698431365
transform -1 0 17248 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2449_
timestamp 1698431365
transform 1 0 12096 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2450_
timestamp 1698431365
transform 1 0 15904 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2451_
timestamp 1698431365
transform 1 0 17248 0 1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2452_
timestamp 1698431365
transform -1 0 21728 0 -1 25088
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2453_
timestamp 1698431365
transform 1 0 38528 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2454_
timestamp 1698431365
transform -1 0 23408 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2455_
timestamp 1698431365
transform -1 0 24864 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2456_
timestamp 1698431365
transform 1 0 10080 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _2457_
timestamp 1698431365
transform 1 0 13328 0 -1 12544
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2458_
timestamp 1698431365
transform 1 0 23632 0 -1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2459_
timestamp 1698431365
transform 1 0 25760 0 -1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _2460_
timestamp 1698431365
transform 1 0 10080 0 1 10976
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2461_
timestamp 1698431365
transform 1 0 27552 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2462_
timestamp 1698431365
transform -1 0 17808 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2463_
timestamp 1698431365
transform 1 0 28560 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2464_
timestamp 1698431365
transform -1 0 28112 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2465_
timestamp 1698431365
transform 1 0 8512 0 1 14112
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2466_
timestamp 1698431365
transform 1 0 6496 0 -1 15680
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_4  _2467_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10752 0 -1 14112
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2468_
timestamp 1698431365
transform 1 0 29456 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _2469_
timestamp 1698431365
transform 1 0 28224 0 -1 17248
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2470_
timestamp 1698431365
transform 1 0 37520 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2471_
timestamp 1698431365
transform 1 0 37744 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2472_
timestamp 1698431365
transform 1 0 38640 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2473_
timestamp 1698431365
transform -1 0 34384 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2474_
timestamp 1698431365
transform -1 0 39088 0 1 18816
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2475_
timestamp 1698431365
transform -1 0 35504 0 1 20384
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2476_
timestamp 1698431365
transform -1 0 31808 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2477_
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2478_
timestamp 1698431365
transform 1 0 30240 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2479_
timestamp 1698431365
transform 1 0 35728 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2480_
timestamp 1698431365
transform 1 0 38640 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2481_
timestamp 1698431365
transform -1 0 39872 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2482_
timestamp 1698431365
transform -1 0 40992 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2483_
timestamp 1698431365
transform -1 0 46592 0 -1 20384
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2484_
timestamp 1698431365
transform 1 0 39872 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2485_
timestamp 1698431365
transform 1 0 39760 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2486_
timestamp 1698431365
transform -1 0 40544 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2487_
timestamp 1698431365
transform 1 0 38528 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2488_
timestamp 1698431365
transform 1 0 41552 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2489_
timestamp 1698431365
transform -1 0 44576 0 -1 20384
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2490_
timestamp 1698431365
transform 1 0 46256 0 1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2491_
timestamp 1698431365
transform 1 0 46256 0 1 20384
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2492_
timestamp 1698431365
transform 1 0 49280 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2493_
timestamp 1698431365
transform 1 0 50624 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _2494_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 46592 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2495_
timestamp 1698431365
transform 1 0 48832 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2496_
timestamp 1698431365
transform -1 0 23296 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2497_
timestamp 1698431365
transform -1 0 26208 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2498_
timestamp 1698431365
transform -1 0 19376 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2499_
timestamp 1698431365
transform 1 0 23856 0 1 15680
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2500_
timestamp 1698431365
transform -1 0 23968 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2501_
timestamp 1698431365
transform -1 0 13664 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _2502_
timestamp 1698431365
transform 1 0 10080 0 1 15680
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2503_
timestamp 1698431365
transform 1 0 10080 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _2504_
timestamp 1698431365
transform -1 0 15680 0 -1 7840
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _2505_
timestamp 1698431365
transform -1 0 22288 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _2506_
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2507_
timestamp 1698431365
transform 1 0 21392 0 -1 14112
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _2508_
timestamp 1698431365
transform 1 0 21504 0 1 12544
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2509_
timestamp 1698431365
transform 1 0 41440 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2510_
timestamp 1698431365
transform -1 0 42112 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2511_
timestamp 1698431365
transform 1 0 42112 0 -1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2512_
timestamp 1698431365
transform 1 0 33040 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2513_
timestamp 1698431365
transform 1 0 35616 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2514_
timestamp 1698431365
transform 1 0 8624 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2515_
timestamp 1698431365
transform 1 0 11088 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2516_
timestamp 1698431365
transform 1 0 11200 0 1 14112
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2517_
timestamp 1698431365
transform -1 0 17472 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2518_
timestamp 1698431365
transform 1 0 14336 0 1 15680
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2519_
timestamp 1698431365
transform -1 0 16464 0 -1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2520_
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2521_
timestamp 1698431365
transform 1 0 7168 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2522_
timestamp 1698431365
transform -1 0 9744 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2523_
timestamp 1698431365
transform 1 0 9744 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2524_
timestamp 1698431365
transform 1 0 11536 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2525_
timestamp 1698431365
transform -1 0 14784 0 -1 10976
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2526_
timestamp 1698431365
transform 1 0 15456 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _2527_
timestamp 1698431365
transform -1 0 16912 0 1 12544
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _2528_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12208 0 -1 15680
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2529_
timestamp 1698431365
transform 1 0 31248 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _2530_
timestamp 1698431365
transform 1 0 31696 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2531_
timestamp 1698431365
transform 1 0 34720 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2532_
timestamp 1698431365
transform -1 0 34048 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2533_
timestamp 1698431365
transform 1 0 30800 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2534_
timestamp 1698431365
transform -1 0 33824 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2535_
timestamp 1698431365
transform -1 0 35616 0 1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _2536_
timestamp 1698431365
transform -1 0 20944 0 1 17248
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2537_
timestamp 1698431365
transform -1 0 21728 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _2538_
timestamp 1698431365
transform -1 0 24864 0 -1 17248
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2539_
timestamp 1698431365
transform -1 0 17920 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2540_
timestamp 1698431365
transform 1 0 22512 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2541_
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _2542_
timestamp 1698431365
transform 1 0 23968 0 1 17248
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2543_
timestamp 1698431365
transform 1 0 38304 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2544_
timestamp 1698431365
transform -1 0 38752 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2545_
timestamp 1698431365
transform 1 0 38976 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2546_
timestamp 1698431365
transform 1 0 45248 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2547_
timestamp 1698431365
transform 1 0 46704 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2548_
timestamp 1698431365
transform 1 0 48944 0 1 17248
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2549_
timestamp 1698431365
transform 1 0 43232 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2550_
timestamp 1698431365
transform 1 0 41552 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2551_
timestamp 1698431365
transform 1 0 40992 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2552_
timestamp 1698431365
transform -1 0 44240 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2553_
timestamp 1698431365
transform 1 0 43904 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2554_
timestamp 1698431365
transform -1 0 44464 0 1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2555_
timestamp 1698431365
transform 1 0 45472 0 1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2556_
timestamp 1698431365
transform 1 0 48832 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2557_
timestamp 1698431365
transform 1 0 49728 0 1 18816
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2558_
timestamp 1698431365
transform 1 0 52528 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2559_
timestamp 1698431365
transform -1 0 47712 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _2560_
timestamp 1698431365
transform -1 0 47376 0 -1 17248
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2561_
timestamp 1698431365
transform -1 0 19264 0 1 12544
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2562_
timestamp 1698431365
transform 1 0 17696 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2563_
timestamp 1698431365
transform 1 0 18816 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2564_
timestamp 1698431365
transform 1 0 18032 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2565_
timestamp 1698431365
transform -1 0 18368 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2566_
timestamp 1698431365
transform 1 0 15792 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _2567_
timestamp 1698431365
transform 1 0 16464 0 1 7840
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _2568_
timestamp 1698431365
transform 1 0 17696 0 -1 12544
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2569_
timestamp 1698431365
transform -1 0 42784 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2570_
timestamp 1698431365
transform -1 0 42336 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2571_
timestamp 1698431365
transform 1 0 42336 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2572_
timestamp 1698431365
transform 1 0 16128 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2573_
timestamp 1698431365
transform 1 0 27552 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2574_
timestamp 1698431365
transform 1 0 9632 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2575_
timestamp 1698431365
transform 1 0 10976 0 -1 12544
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2576_
timestamp 1698431365
transform 1 0 24304 0 1 14112
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2577_
timestamp 1698431365
transform 1 0 20832 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2578_
timestamp 1698431365
transform -1 0 27888 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2579_
timestamp 1698431365
transform 1 0 30128 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2580_
timestamp 1698431365
transform -1 0 35504 0 -1 14112
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2581_
timestamp 1698431365
transform -1 0 34720 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2582_
timestamp 1698431365
transform -1 0 32704 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2583_
timestamp 1698431365
transform -1 0 30688 0 1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2584_
timestamp 1698431365
transform -1 0 33824 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2585_
timestamp 1698431365
transform 1 0 41888 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2586_
timestamp 1698431365
transform 1 0 18704 0 -1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2587_
timestamp 1698431365
transform 1 0 19712 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2588_
timestamp 1698431365
transform 1 0 29232 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2589_
timestamp 1698431365
transform 1 0 29008 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2590_
timestamp 1698431365
transform 1 0 29344 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2591_
timestamp 1698431365
transform 1 0 23184 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2592_
timestamp 1698431365
transform 1 0 31920 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2593_
timestamp 1698431365
transform -1 0 36288 0 1 17248
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2594_
timestamp 1698431365
transform 1 0 38304 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2595_
timestamp 1698431365
transform -1 0 37968 0 -1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2596_
timestamp 1698431365
transform 1 0 28112 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2597_
timestamp 1698431365
transform 1 0 28784 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2598_
timestamp 1698431365
transform 1 0 23184 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2599_
timestamp 1698431365
transform -1 0 14560 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2600_
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2601_
timestamp 1698431365
transform 1 0 23296 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2602_
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2603_
timestamp 1698431365
transform -1 0 25200 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _2604_
timestamp 1698431365
transform 1 0 25200 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2605_
timestamp 1698431365
transform -1 0 17136 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2606_
timestamp 1698431365
transform 1 0 12096 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2607_
timestamp 1698431365
transform 1 0 14672 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2608_
timestamp 1698431365
transform -1 0 16016 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2609_
timestamp 1698431365
transform -1 0 15008 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2610_
timestamp 1698431365
transform 1 0 13328 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai33_1  _2611_
timestamp 1698431365
transform 1 0 13664 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2612_
timestamp 1698431365
transform 1 0 27328 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2613_
timestamp 1698431365
transform 1 0 36624 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2614_
timestamp 1698431365
transform -1 0 39648 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2615_
timestamp 1698431365
transform 1 0 44688 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2616_
timestamp 1698431365
transform 1 0 41104 0 1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2617_
timestamp 1698431365
transform 1 0 37072 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2618_
timestamp 1698431365
transform 1 0 37632 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2619_
timestamp 1698431365
transform -1 0 44464 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2620_
timestamp 1698431365
transform 1 0 47152 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2621_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 46816 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2622_
timestamp 1698431365
transform 1 0 49056 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2623_
timestamp 1698431365
transform 1 0 47600 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2624_
timestamp 1698431365
transform -1 0 50960 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2625_
timestamp 1698431365
transform 1 0 50960 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2626_
timestamp 1698431365
transform 1 0 50400 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2627_
timestamp 1698431365
transform 1 0 52528 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2628_
timestamp 1698431365
transform 1 0 45248 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2629_
timestamp 1698431365
transform -1 0 43792 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2630_
timestamp 1698431365
transform 1 0 45696 0 -1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2631_
timestamp 1698431365
transform 1 0 17584 0 -1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2632_
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2633_
timestamp 1698431365
transform 1 0 25424 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2634_
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2635_
timestamp 1698431365
transform -1 0 22848 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2636_
timestamp 1698431365
transform -1 0 21840 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2637_
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2638_
timestamp 1698431365
transform 1 0 26320 0 -1 6272
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2639_
timestamp 1698431365
transform 1 0 27104 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2640_
timestamp 1698431365
transform -1 0 42784 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2641_
timestamp 1698431365
transform 1 0 43568 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2642_
timestamp 1698431365
transform 1 0 42896 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2643_
timestamp 1698431365
transform -1 0 35616 0 1 14112
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2644_
timestamp 1698431365
transform 1 0 26320 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2645_
timestamp 1698431365
transform 1 0 25872 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2646_
timestamp 1698431365
transform 1 0 19712 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2647_
timestamp 1698431365
transform 1 0 21056 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2648_
timestamp 1698431365
transform -1 0 28224 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2649_
timestamp 1698431365
transform 1 0 26432 0 1 15680
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2650_
timestamp 1698431365
transform -1 0 30128 0 -1 14112
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2651_
timestamp 1698431365
transform -1 0 36736 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2652_
timestamp 1698431365
transform 1 0 35616 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2653_
timestamp 1698431365
transform 1 0 33712 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2654_
timestamp 1698431365
transform -1 0 38192 0 -1 17248
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2655_
timestamp 1698431365
transform -1 0 39424 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _2656_
timestamp 1698431365
transform 1 0 37968 0 -1 15680
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2657_
timestamp 1698431365
transform 1 0 39088 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2658_
timestamp 1698431365
transform -1 0 38528 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2659_
timestamp 1698431365
transform 1 0 38976 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2660_
timestamp 1698431365
transform -1 0 41328 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _2661_
timestamp 1698431365
transform 1 0 39536 0 1 15680
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2662_
timestamp 1698431365
transform 1 0 45248 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2663_
timestamp 1698431365
transform 1 0 46256 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2664_
timestamp 1698431365
transform 1 0 49728 0 1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2665_
timestamp 1698431365
transform 1 0 46144 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2666_
timestamp 1698431365
transform -1 0 46032 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2667_
timestamp 1698431365
transform 1 0 44688 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2668_
timestamp 1698431365
transform 1 0 45584 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2669_
timestamp 1698431365
transform -1 0 48384 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2670_
timestamp 1698431365
transform -1 0 50400 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2671_
timestamp 1698431365
transform 1 0 50848 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2672_
timestamp 1698431365
transform 1 0 51408 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2673_
timestamp 1698431365
transform 1 0 52864 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2674_
timestamp 1698431365
transform 1 0 46256 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2675_
timestamp 1698431365
transform 1 0 47152 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2676_
timestamp 1698431365
transform 1 0 42112 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2677_
timestamp 1698431365
transform 1 0 24192 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2678_
timestamp 1698431365
transform 1 0 13664 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2679_
timestamp 1698431365
transform -1 0 21056 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2680_
timestamp 1698431365
transform 1 0 21728 0 -1 25088
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2681_
timestamp 1698431365
transform 1 0 23744 0 -1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2682_
timestamp 1698431365
transform 1 0 26768 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2683_
timestamp 1698431365
transform -1 0 28448 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2684_
timestamp 1698431365
transform 1 0 25984 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _2685_
timestamp 1698431365
transform 1 0 26320 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2686_
timestamp 1698431365
transform 1 0 41888 0 -1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _2687_
timestamp 1698431365
transform 1 0 29792 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2688_
timestamp 1698431365
transform 1 0 31920 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2689_
timestamp 1698431365
transform -1 0 28784 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2690_
timestamp 1698431365
transform 1 0 11424 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2691_
timestamp 1698431365
transform -1 0 22176 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2692_
timestamp 1698431365
transform -1 0 20944 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2693_
timestamp 1698431365
transform -1 0 20048 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2694_
timestamp 1698431365
transform 1 0 18928 0 -1 4704
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2695_
timestamp 1698431365
transform 1 0 21280 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2696_
timestamp 1698431365
transform -1 0 22960 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2697_
timestamp 1698431365
transform 1 0 31360 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2698_
timestamp 1698431365
transform 1 0 18816 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2699_
timestamp 1698431365
transform 1 0 19264 0 1 6272
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2700_
timestamp 1698431365
transform -1 0 20944 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2701_
timestamp 1698431365
transform 1 0 17472 0 1 4704
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2702_
timestamp 1698431365
transform 1 0 22064 0 -1 4704
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2703_
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2704_
timestamp 1698431365
transform 1 0 22512 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2705_
timestamp 1698431365
transform 1 0 21840 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2706_
timestamp 1698431365
transform 1 0 38304 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2707_
timestamp 1698431365
transform 1 0 38864 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2708_
timestamp 1698431365
transform 1 0 44352 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2709_
timestamp 1698431365
transform -1 0 44464 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2710_
timestamp 1698431365
transform -1 0 46368 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2711_
timestamp 1698431365
transform 1 0 46368 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _2712_
timestamp 1698431365
transform 1 0 48608 0 -1 10976
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2713_
timestamp 1698431365
transform 1 0 49840 0 -1 17248
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2714_
timestamp 1698431365
transform 1 0 48832 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2715_
timestamp 1698431365
transform 1 0 49952 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2716_
timestamp 1698431365
transform 1 0 51520 0 -1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2717_
timestamp 1698431365
transform 1 0 48832 0 -1 14112
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2718_
timestamp 1698431365
transform 1 0 49840 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2719_
timestamp 1698431365
transform 1 0 51184 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2720_
timestamp 1698431365
transform 1 0 46368 0 1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2721_
timestamp 1698431365
transform -1 0 42224 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2722_
timestamp 1698431365
transform -1 0 16016 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _2723_
timestamp 1698431365
transform 1 0 16016 0 1 6272
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2724_
timestamp 1698431365
transform -1 0 17024 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2725_
timestamp 1698431365
transform 1 0 23968 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2726_
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2727_
timestamp 1698431365
transform 1 0 31248 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2728_
timestamp 1698431365
transform -1 0 36288 0 -1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2729_
timestamp 1698431365
transform -1 0 15680 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2730_
timestamp 1698431365
transform -1 0 24640 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2731_
timestamp 1698431365
transform -1 0 16128 0 -1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2732_
timestamp 1698431365
transform -1 0 12208 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2733_
timestamp 1698431365
transform -1 0 16352 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _2734_
timestamp 1698431365
transform -1 0 18816 0 1 10976
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2735_
timestamp 1698431365
transform 1 0 33040 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2736_
timestamp 1698431365
transform 1 0 33040 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2737_
timestamp 1698431365
transform 1 0 40208 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2738_
timestamp 1698431365
transform -1 0 43344 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2739_
timestamp 1698431365
transform 1 0 42224 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2740_
timestamp 1698431365
transform -1 0 46256 0 1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2741_
timestamp 1698431365
transform -1 0 36064 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2742_
timestamp 1698431365
transform 1 0 25312 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2743_
timestamp 1698431365
transform -1 0 28784 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2744_
timestamp 1698431365
transform 1 0 19040 0 1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2745_
timestamp 1698431365
transform 1 0 18368 0 -1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2746_
timestamp 1698431365
transform 1 0 24304 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2747_
timestamp 1698431365
transform 1 0 25312 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2748_
timestamp 1698431365
transform 1 0 34944 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2749_
timestamp 1698431365
transform 1 0 45248 0 -1 7840
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _2750_
timestamp 1698431365
transform 1 0 47488 0 1 6272
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2751_
timestamp 1698431365
transform 1 0 48832 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2752_
timestamp 1698431365
transform 1 0 50400 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2753_
timestamp 1698431365
transform 1 0 51072 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2754_
timestamp 1698431365
transform 1 0 50176 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2755_
timestamp 1698431365
transform 1 0 51520 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2756_
timestamp 1698431365
transform -1 0 46368 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2757_
timestamp 1698431365
transform 1 0 22400 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2758_
timestamp 1698431365
transform 1 0 23632 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2759_
timestamp 1698431365
transform 1 0 23408 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2760_
timestamp 1698431365
transform 1 0 24752 0 1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2761_
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2762_
timestamp 1698431365
transform -1 0 40768 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2763_
timestamp 1698431365
transform 1 0 33264 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2764_
timestamp 1698431365
transform 1 0 24528 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2765_
timestamp 1698431365
transform 1 0 29680 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2766_
timestamp 1698431365
transform -1 0 29120 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2767_
timestamp 1698431365
transform -1 0 27216 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2768_
timestamp 1698431365
transform -1 0 30464 0 1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2769_
timestamp 1698431365
transform 1 0 31248 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2770_
timestamp 1698431365
transform 1 0 31360 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2771_
timestamp 1698431365
transform -1 0 33600 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2772_
timestamp 1698431365
transform -1 0 33488 0 1 3136
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2773_
timestamp 1698431365
transform -1 0 42000 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _2774_
timestamp 1698431365
transform 1 0 19152 0 -1 9408
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2775_
timestamp 1698431365
transform 1 0 29792 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2776_
timestamp 1698431365
transform 1 0 30688 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2777_
timestamp 1698431365
transform 1 0 31024 0 -1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2778_
timestamp 1698431365
transform 1 0 46144 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2779_
timestamp 1698431365
transform -1 0 50400 0 -1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2780_
timestamp 1698431365
transform -1 0 49952 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _2781_
timestamp 1698431365
transform -1 0 51520 0 1 7840
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2782_
timestamp 1698431365
transform 1 0 49168 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2783_
timestamp 1698431365
transform 1 0 50512 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2784_
timestamp 1698431365
transform -1 0 33824 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2785_
timestamp 1698431365
transform -1 0 31024 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2786_
timestamp 1698431365
transform 1 0 45024 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2787_
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2788_
timestamp 1698431365
transform 1 0 29456 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2789_
timestamp 1698431365
transform 1 0 30464 0 -1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2790_
timestamp 1698431365
transform 1 0 34720 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2791_
timestamp 1698431365
transform 1 0 17696 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2792_
timestamp 1698431365
transform 1 0 20384 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2793_
timestamp 1698431365
transform -1 0 25200 0 1 21952
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2794_
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2795_
timestamp 1698431365
transform 1 0 34160 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2796_
timestamp 1698431365
transform 1 0 34720 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2797_
timestamp 1698431365
transform 1 0 34608 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2798_
timestamp 1698431365
transform -1 0 29904 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2799_
timestamp 1698431365
transform 1 0 27440 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2800_
timestamp 1698431365
transform 1 0 28112 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2801_
timestamp 1698431365
transform 1 0 29904 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2802_
timestamp 1698431365
transform 1 0 32928 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2803_
timestamp 1698431365
transform 1 0 33264 0 -1 7840
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2804_
timestamp 1698431365
transform 1 0 34384 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2805_
timestamp 1698431365
transform 1 0 33824 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2806_
timestamp 1698431365
transform -1 0 35840 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2807_
timestamp 1698431365
transform 1 0 34720 0 -1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2808_
timestamp 1698431365
transform 1 0 47488 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2809_
timestamp 1698431365
transform 1 0 48608 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2810_
timestamp 1698431365
transform -1 0 51520 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2811_
timestamp 1698431365
transform 1 0 48608 0 -1 4704
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2812_
timestamp 1698431365
transform 1 0 50288 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2813_
timestamp 1698431365
transform -1 0 22064 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2814_
timestamp 1698431365
transform -1 0 27888 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2815_
timestamp 1698431365
transform 1 0 38304 0 -1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2816_
timestamp 1698431365
transform 1 0 38080 0 -1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2817_
timestamp 1698431365
transform 1 0 39536 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2818_
timestamp 1698431365
transform -1 0 30128 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2819_
timestamp 1698431365
transform -1 0 35840 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2820_
timestamp 1698431365
transform 1 0 32480 0 1 6272
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2821_
timestamp 1698431365
transform -1 0 39536 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2822_
timestamp 1698431365
transform -1 0 36624 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2823_
timestamp 1698431365
transform -1 0 37632 0 -1 12544
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2824_
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2825_
timestamp 1698431365
transform 1 0 37744 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2826_
timestamp 1698431365
transform -1 0 34720 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2827_
timestamp 1698431365
transform 1 0 37856 0 -1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2828_
timestamp 1698431365
transform -1 0 47600 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2829_
timestamp 1698431365
transform 1 0 49280 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2830_
timestamp 1698431365
transform -1 0 49280 0 1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2831_
timestamp 1698431365
transform -1 0 46928 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2832_
timestamp 1698431365
transform 1 0 44912 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2833_
timestamp 1698431365
transform 1 0 46928 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2834_
timestamp 1698431365
transform 1 0 39536 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2835_
timestamp 1698431365
transform 1 0 39200 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2836_
timestamp 1698431365
transform -1 0 20944 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2837_
timestamp 1698431365
transform 1 0 23072 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2838_
timestamp 1698431365
transform 1 0 23968 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2839_
timestamp 1698431365
transform 1 0 35840 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2840_
timestamp 1698431365
transform -1 0 37744 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2841_
timestamp 1698431365
transform 1 0 37744 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2842_
timestamp 1698431365
transform -1 0 38080 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2843_
timestamp 1698431365
transform 1 0 35280 0 -1 6272
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2844_
timestamp 1698431365
transform -1 0 41664 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2845_
timestamp 1698431365
transform 1 0 40208 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2846_
timestamp 1698431365
transform 1 0 41440 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2847_
timestamp 1698431365
transform 1 0 42672 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2848_
timestamp 1698431365
transform 1 0 38416 0 1 3136
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2849_
timestamp 1698431365
transform 1 0 42784 0 -1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2850_
timestamp 1698431365
transform 1 0 42560 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2851_
timestamp 1698431365
transform 1 0 43120 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2852_
timestamp 1698431365
transform 1 0 38864 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2853_
timestamp 1698431365
transform -1 0 38864 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2854_
timestamp 1698431365
transform 1 0 38528 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2855_
timestamp 1698431365
transform 1 0 43904 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2856_
timestamp 1698431365
transform 1 0 44016 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2857_
timestamp 1698431365
transform 1 0 39312 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2858_
timestamp 1698431365
transform -1 0 42560 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _2859_
timestamp 1698431365
transform 1 0 41664 0 -1 7840
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2860_
timestamp 1698431365
transform 1 0 48608 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2861_
timestamp 1698431365
transform 1 0 49616 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2862_
timestamp 1698431365
transform 1 0 33152 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2863_
timestamp 1698431365
transform 1 0 32816 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2864_
timestamp 1698431365
transform 1 0 31472 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2865_
timestamp 1698431365
transform -1 0 31248 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2866_
timestamp 1698431365
transform 1 0 26320 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2867_
timestamp 1698431365
transform 1 0 25312 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2868_
timestamp 1698431365
transform -1 0 34048 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2869_
timestamp 1698431365
transform 1 0 33712 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2870_
timestamp 1698431365
transform 1 0 17360 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2871_
timestamp 1698431365
transform -1 0 11312 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2872_
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2873_
timestamp 1698431365
transform 1 0 18816 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2874_
timestamp 1698431365
transform 1 0 17696 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2875_
timestamp 1698431365
transform 1 0 18256 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2876_
timestamp 1698431365
transform -1 0 18704 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2877_
timestamp 1698431365
transform -1 0 18144 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2878_
timestamp 1698431365
transform -1 0 6160 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2879_
timestamp 1698431365
transform 1 0 19600 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2880_
timestamp 1698431365
transform -1 0 20608 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2881_
timestamp 1698431365
transform 1 0 13440 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2882_
timestamp 1698431365
transform 1 0 22064 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2883_
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2884_
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2885_
timestamp 1698431365
transform -1 0 22064 0 -1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2886_
timestamp 1698431365
transform 1 0 18032 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2887_
timestamp 1698431365
transform 1 0 23296 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2888_
timestamp 1698431365
transform 1 0 23632 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2889_
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2890_
timestamp 1698431365
transform -1 0 20160 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2891_
timestamp 1698431365
transform 1 0 19936 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2892_
timestamp 1698431365
transform -1 0 23296 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2893_
timestamp 1698431365
transform 1 0 21840 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2894_
timestamp 1698431365
transform -1 0 20384 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2895_
timestamp 1698431365
transform 1 0 20720 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2896_
timestamp 1698431365
transform -1 0 19936 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2897_
timestamp 1698431365
transform -1 0 25872 0 -1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2898_
timestamp 1698431365
transform -1 0 27216 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2899_
timestamp 1698431365
transform -1 0 26544 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2900_
timestamp 1698431365
transform -1 0 25424 0 1 32928
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2901_
timestamp 1698431365
transform 1 0 25424 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2902_
timestamp 1698431365
transform -1 0 26656 0 1 32928
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2903_
timestamp 1698431365
transform -1 0 46144 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2904_
timestamp 1698431365
transform -1 0 44464 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2905_
timestamp 1698431365
transform -1 0 32256 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2906_
timestamp 1698431365
transform 1 0 30800 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2907_
timestamp 1698431365
transform -1 0 29680 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2908_
timestamp 1698431365
transform -1 0 43680 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2909_
timestamp 1698431365
transform -1 0 43120 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2910_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33152 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2911_
timestamp 1698431365
transform 1 0 29792 0 1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2912_
timestamp 1698431365
transform 1 0 33488 0 -1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2913_
timestamp 1698431365
transform -1 0 11536 0 1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2914_
timestamp 1698431365
transform 1 0 4368 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2915_
timestamp 1698431365
transform 1 0 4704 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2916_
timestamp 1698431365
transform -1 0 16240 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  _2917_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 25200 0 1 31360
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  _2918_
timestamp 1698431365
transform 1 0 24752 0 1 29792
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2919_
timestamp 1698431365
transform -1 0 12320 0 1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2920_
timestamp 1698431365
transform 1 0 5376 0 -1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2921_
timestamp 1698431365
transform -1 0 9296 0 1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2922_
timestamp 1698431365
transform -1 0 14336 0 -1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  _2923_
timestamp 1698431365
transform -1 0 17808 0 1 32928
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2924_
timestamp 1698431365
transform 1 0 26096 0 -1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2925_
timestamp 1698431365
transform 1 0 42672 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2926_
timestamp 1698431365
transform 1 0 42448 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _2927_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 35840 0 -1 28224
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2928_
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2929_
timestamp 1698431365
transform 1 0 31024 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2930_
timestamp 1698431365
transform 1 0 27888 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _2931_
timestamp 1698431365
transform 1 0 39760 0 1 29792
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2932_
timestamp 1698431365
transform -1 0 41216 0 1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2933_
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2934_
timestamp 1698431365
transform 1 0 42224 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2935_
timestamp 1698431365
transform 1 0 38528 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1455__A1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1456__I
timestamp 1698431365
transform 1 0 24640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1457__A1
timestamp 1698431365
transform 1 0 29008 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1468__I
timestamp 1698431365
transform 1 0 26880 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1469__I
timestamp 1698431365
transform 1 0 29792 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1470__A1
timestamp 1698431365
transform 1 0 22736 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1474__A2
timestamp 1698431365
transform 1 0 24192 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1475__I
timestamp 1698431365
transform 1 0 27664 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1477__A1
timestamp 1698431365
transform -1 0 21616 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1478__A2
timestamp 1698431365
transform 1 0 29680 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1478__B
timestamp 1698431365
transform 1 0 30688 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1478__C
timestamp 1698431365
transform -1 0 28560 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1479__A1
timestamp 1698431365
transform 1 0 31248 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1487__I
timestamp 1698431365
transform -1 0 10976 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1488__I
timestamp 1698431365
transform 1 0 12880 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1494__A1
timestamp 1698431365
transform 1 0 21168 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1497__I
timestamp 1698431365
transform -1 0 8848 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1500__I
timestamp 1698431365
transform -1 0 8176 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1504__A1
timestamp 1698431365
transform -1 0 24080 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1504__A2
timestamp 1698431365
transform -1 0 23632 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1506__I
timestamp 1698431365
transform 1 0 11872 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1508__A2
timestamp 1698431365
transform -1 0 16576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1509__B
timestamp 1698431365
transform 1 0 25984 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1513__I
timestamp 1698431365
transform 1 0 12432 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1520__A1
timestamp 1698431365
transform 1 0 29792 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1520__A2
timestamp 1698431365
transform 1 0 27440 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1520__B
timestamp 1698431365
transform 1 0 33152 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1521__A1
timestamp 1698431365
transform 1 0 33824 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1521__A3
timestamp 1698431365
transform 1 0 33376 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1523__I
timestamp 1698431365
transform 1 0 32032 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1531__A1
timestamp 1698431365
transform 1 0 37856 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1534__I
timestamp 1698431365
transform 1 0 38416 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1545__I
timestamp 1698431365
transform 1 0 35392 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1558__I
timestamp 1698431365
transform 1 0 17472 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1559__A2
timestamp 1698431365
transform 1 0 25984 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1564__I
timestamp 1698431365
transform 1 0 8400 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1567__I
timestamp 1698431365
transform 1 0 29344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1571__A1
timestamp 1698431365
transform 1 0 16800 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1571__B
timestamp 1698431365
transform 1 0 22064 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1575__B2
timestamp 1698431365
transform 1 0 32368 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1581__I
timestamp 1698431365
transform 1 0 23296 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1584__I
timestamp 1698431365
transform 1 0 19152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1587__A2
timestamp 1698431365
transform 1 0 23072 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1587__B
timestamp 1698431365
transform 1 0 23520 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1588__A2
timestamp 1698431365
transform -1 0 18928 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1588__B
timestamp 1698431365
transform -1 0 17248 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1589__A1
timestamp 1698431365
transform 1 0 35952 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1590__A1
timestamp 1698431365
transform 1 0 46144 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1591__I
timestamp 1698431365
transform 1 0 46928 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1594__I
timestamp 1698431365
transform 1 0 16800 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1595__I
timestamp 1698431365
transform -1 0 16128 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1601__A2
timestamp 1698431365
transform 1 0 10528 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1605__A1
timestamp 1698431365
transform 1 0 11760 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1606__A2
timestamp 1698431365
transform 1 0 29232 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1607__A3
timestamp 1698431365
transform -1 0 12992 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1607__B
timestamp 1698431365
transform -1 0 15680 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1611__A1
timestamp 1698431365
transform 1 0 15680 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1611__B
timestamp 1698431365
transform -1 0 18368 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1612__I
timestamp 1698431365
transform 1 0 8624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1615__A3
timestamp 1698431365
transform -1 0 9296 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1617__A1
timestamp 1698431365
transform 1 0 12880 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1618__A1
timestamp 1698431365
transform -1 0 11424 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1619__I0
timestamp 1698431365
transform -1 0 11424 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1620__I
timestamp 1698431365
transform -1 0 13888 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1622__I
timestamp 1698431365
transform -1 0 47824 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1625__I
timestamp 1698431365
transform 1 0 11088 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1627__I
timestamp 1698431365
transform -1 0 15232 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1636__A2
timestamp 1698431365
transform 1 0 20720 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1642__A1
timestamp 1698431365
transform -1 0 13888 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1642__B
timestamp 1698431365
transform 1 0 12432 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1643__A1
timestamp 1698431365
transform -1 0 13440 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1645__A1
timestamp 1698431365
transform 1 0 23744 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1645__B1
timestamp 1698431365
transform 1 0 15232 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1646__A1
timestamp 1698431365
transform 1 0 37968 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1646__A2
timestamp 1698431365
transform 1 0 38416 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1648__A1
timestamp 1698431365
transform 1 0 38976 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1649__A1
timestamp 1698431365
transform 1 0 41776 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1654__I
timestamp 1698431365
transform 1 0 36960 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1655__I
timestamp 1698431365
transform 1 0 34832 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1656__I
timestamp 1698431365
transform 1 0 36512 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1657__I
timestamp 1698431365
transform -1 0 17696 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1658__A3
timestamp 1698431365
transform 1 0 19376 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1659__A2
timestamp 1698431365
transform 1 0 37408 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1660__A2
timestamp 1698431365
transform -1 0 26880 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1660__B1
timestamp 1698431365
transform 1 0 36400 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1663__A1
timestamp 1698431365
transform -1 0 23968 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1663__B
timestamp 1698431365
transform -1 0 25648 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1665__I
timestamp 1698431365
transform 1 0 18256 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__A2
timestamp 1698431365
transform -1 0 26656 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1667__A1
timestamp 1698431365
transform 1 0 14112 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1669__A1
timestamp 1698431365
transform -1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1669__A2
timestamp 1698431365
transform 1 0 11984 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1672__A1
timestamp 1698431365
transform 1 0 34048 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1672__C2
timestamp 1698431365
transform 1 0 33152 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1673__A1
timestamp 1698431365
transform -1 0 44576 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1675__A1
timestamp 1698431365
transform 1 0 39088 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1676__I
timestamp 1698431365
transform 1 0 18816 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1678__A2
timestamp 1698431365
transform -1 0 10864 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1679__A1
timestamp 1698431365
transform 1 0 22288 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1683__A1
timestamp 1698431365
transform 1 0 20496 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1688__I1
timestamp 1698431365
transform 1 0 16352 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1688__S0
timestamp 1698431365
transform 1 0 16800 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1690__A1
timestamp 1698431365
transform 1 0 31472 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1693__I
timestamp 1698431365
transform 1 0 18256 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1695__A1
timestamp 1698431365
transform -1 0 18032 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1695__A2
timestamp 1698431365
transform -1 0 17584 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1695__B
timestamp 1698431365
transform -1 0 16352 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1697__A1
timestamp 1698431365
transform 1 0 18032 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1698__C
timestamp 1698431365
transform -1 0 18144 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1701__A2
timestamp 1698431365
transform -1 0 10416 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1702__B
timestamp 1698431365
transform -1 0 10080 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1705__A1
timestamp 1698431365
transform -1 0 12544 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1705__C
timestamp 1698431365
transform -1 0 14000 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1706__A2
timestamp 1698431365
transform -1 0 13440 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1707__A1
timestamp 1698431365
transform -1 0 21168 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1710__I
timestamp 1698431365
transform 1 0 46704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1714__B
timestamp 1698431365
transform 1 0 13552 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1718__A3
timestamp 1698431365
transform -1 0 13776 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1721__A1
timestamp 1698431365
transform 1 0 29456 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1721__A2
timestamp 1698431365
transform 1 0 33264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1722__A1
timestamp 1698431365
transform -1 0 29680 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1722__A2
timestamp 1698431365
transform 1 0 27552 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1723__A1
timestamp 1698431365
transform 1 0 34496 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1725__A2
timestamp 1698431365
transform -1 0 39760 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1725__A3
timestamp 1698431365
transform -1 0 39312 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1727__I
timestamp 1698431365
transform 1 0 38976 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1728__I
timestamp 1698431365
transform 1 0 18816 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1735__I
timestamp 1698431365
transform 1 0 17696 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1736__A2
timestamp 1698431365
transform -1 0 21504 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1736__A3
timestamp 1698431365
transform 1 0 21504 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1737__A2
timestamp 1698431365
transform -1 0 22848 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1741__A1
timestamp 1698431365
transform 1 0 27328 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1743__B
timestamp 1698431365
transform 1 0 26208 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1746__A1
timestamp 1698431365
transform 1 0 33152 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1746__A2
timestamp 1698431365
transform -1 0 30464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1747__A2
timestamp 1698431365
transform -1 0 16800 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1749__A2
timestamp 1698431365
transform 1 0 33712 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1749__B
timestamp 1698431365
transform -1 0 26992 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1761__A1
timestamp 1698431365
transform 1 0 33600 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1763__A1
timestamp 1698431365
transform -1 0 38864 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1765__A2
timestamp 1698431365
transform 1 0 26544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1766__I
timestamp 1698431365
transform -1 0 13888 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1767__A1
timestamp 1698431365
transform -1 0 18592 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1772__A2
timestamp 1698431365
transform 1 0 23408 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1775__A2
timestamp 1698431365
transform 1 0 19488 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1779__A1
timestamp 1698431365
transform 1 0 23856 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1784__I
timestamp 1698431365
transform -1 0 46816 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1785__I
timestamp 1698431365
transform 1 0 41664 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1786__C
timestamp 1698431365
transform 1 0 34944 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1793__A1
timestamp 1698431365
transform -1 0 7728 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1793__A2
timestamp 1698431365
transform -1 0 10752 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1795__A1
timestamp 1698431365
transform -1 0 13216 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1796__A2
timestamp 1698431365
transform 1 0 20048 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1796__B
timestamp 1698431365
transform 1 0 17920 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1797__A1
timestamp 1698431365
transform -1 0 30352 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1798__B
timestamp 1698431365
transform 1 0 19040 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1799__A2
timestamp 1698431365
transform -1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1800__A1
timestamp 1698431365
transform 1 0 36400 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1805__A1
timestamp 1698431365
transform 1 0 40096 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1805__A2
timestamp 1698431365
transform 1 0 38864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1808__A2
timestamp 1698431365
transform -1 0 14784 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1813__A1
timestamp 1698431365
transform -1 0 23520 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1818__B1
timestamp 1698431365
transform -1 0 16128 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1820__A1
timestamp 1698431365
transform -1 0 24192 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1831__B
timestamp 1698431365
transform 1 0 37968 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1835__A2
timestamp 1698431365
transform -1 0 26544 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1837__A1
timestamp 1698431365
transform 1 0 25424 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1837__A2
timestamp 1698431365
transform 1 0 31024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1838__A2
timestamp 1698431365
transform -1 0 27104 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1839__A1
timestamp 1698431365
transform 1 0 24192 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1840__A1
timestamp 1698431365
transform 1 0 24640 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1841__B2
timestamp 1698431365
transform 1 0 30240 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1843__A2
timestamp 1698431365
transform -1 0 31360 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1843__B
timestamp 1698431365
transform 1 0 30688 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1844__B
timestamp 1698431365
transform 1 0 32032 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1852__A1
timestamp 1698431365
transform 1 0 12432 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1852__A2
timestamp 1698431365
transform -1 0 12096 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1854__A2
timestamp 1698431365
transform -1 0 11760 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1855__A2
timestamp 1698431365
transform 1 0 14000 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1857__A3
timestamp 1698431365
transform -1 0 15008 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1860__C
timestamp 1698431365
transform 1 0 15680 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1862__B2
timestamp 1698431365
transform 1 0 16352 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1864__A1
timestamp 1698431365
transform 1 0 42112 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1866__A1
timestamp 1698431365
transform 1 0 19712 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1870__A1
timestamp 1698431365
transform -1 0 14112 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1870__A2
timestamp 1698431365
transform 1 0 15232 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1871__A1
timestamp 1698431365
transform -1 0 18816 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1872__A2
timestamp 1698431365
transform -1 0 13664 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1873__C
timestamp 1698431365
transform -1 0 21840 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1874__A1
timestamp 1698431365
transform -1 0 40544 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1874__A3
timestamp 1698431365
transform -1 0 38080 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1879__A1
timestamp 1698431365
transform 1 0 48048 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1883__I
timestamp 1698431365
transform -1 0 47264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1884__A1
timestamp 1698431365
transform -1 0 47488 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1892__A1
timestamp 1698431365
transform 1 0 25872 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1892__A2
timestamp 1698431365
transform 1 0 26320 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1897__B2
timestamp 1698431365
transform -1 0 24304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1897__C
timestamp 1698431365
transform 1 0 25984 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1898__I
timestamp 1698431365
transform 1 0 30240 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1899__I
timestamp 1698431365
transform -1 0 27216 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1901__A1
timestamp 1698431365
transform -1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1907__A1
timestamp 1698431365
transform 1 0 38976 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1910__A3
timestamp 1698431365
transform 1 0 47152 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1911__A1
timestamp 1698431365
transform 1 0 11984 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1914__A1
timestamp 1698431365
transform 1 0 12880 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1917__A1
timestamp 1698431365
transform -1 0 20384 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1918__I
timestamp 1698431365
transform -1 0 44912 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1921__A1
timestamp 1698431365
transform 1 0 39424 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1921__A4
timestamp 1698431365
transform 1 0 38976 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1923__B
timestamp 1698431365
transform -1 0 22400 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1925__A2
timestamp 1698431365
transform 1 0 25760 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1927__A1
timestamp 1698431365
transform 1 0 22736 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1928__A2
timestamp 1698431365
transform -1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1931__A1
timestamp 1698431365
transform 1 0 27664 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1932__A2
timestamp 1698431365
transform -1 0 38416 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1946__A1
timestamp 1698431365
transform 1 0 49616 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1950__I
timestamp 1698431365
transform 1 0 30352 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1951__A3
timestamp 1698431365
transform 1 0 28560 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1952__B
timestamp 1698431365
transform 1 0 25312 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1955__A1
timestamp 1698431365
transform -1 0 31472 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1959__A3
timestamp 1698431365
transform 1 0 40992 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1959__A4
timestamp 1698431365
transform 1 0 41440 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1960__A2
timestamp 1698431365
transform 1 0 19824 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1960__B
timestamp 1698431365
transform -1 0 18816 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1963__A2
timestamp 1698431365
transform 1 0 19040 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1965__A1
timestamp 1698431365
transform 1 0 36288 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1970__A1
timestamp 1698431365
transform 1 0 37072 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1970__A4
timestamp 1698431365
transform -1 0 37296 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1972__A2
timestamp 1698431365
transform 1 0 27664 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1975__A2
timestamp 1698431365
transform -1 0 23184 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1975__A3
timestamp 1698431365
transform 1 0 23408 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1976__A1
timestamp 1698431365
transform -1 0 23072 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1976__A2
timestamp 1698431365
transform 1 0 20944 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1977__A2
timestamp 1698431365
transform -1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1977__B
timestamp 1698431365
transform 1 0 33376 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1978__A1
timestamp 1698431365
transform 1 0 33152 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1978__A3
timestamp 1698431365
transform 1 0 32816 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1979__A1
timestamp 1698431365
transform -1 0 34832 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1980__C
timestamp 1698431365
transform 1 0 37968 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1983__A1
timestamp 1698431365
transform 1 0 34608 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2001__I
timestamp 1698431365
transform -1 0 22512 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2002__B
timestamp 1698431365
transform 1 0 24192 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2006__A2
timestamp 1698431365
transform 1 0 34160 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2007__A1
timestamp 1698431365
transform -1 0 33824 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2007__A2
timestamp 1698431365
transform -1 0 34272 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2012__A1
timestamp 1698431365
transform 1 0 26992 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2013__A2
timestamp 1698431365
transform -1 0 29792 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2017__A2
timestamp 1698431365
transform 1 0 28784 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2018__A1
timestamp 1698431365
transform 1 0 30128 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2018__B2
timestamp 1698431365
transform 1 0 25984 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2019__A2
timestamp 1698431365
transform 1 0 44464 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2021__A1
timestamp 1698431365
transform 1 0 34272 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2021__A2
timestamp 1698431365
transform 1 0 33824 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2022__A1
timestamp 1698431365
transform -1 0 33488 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2022__A2
timestamp 1698431365
transform 1 0 33712 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2024__A1
timestamp 1698431365
transform 1 0 22960 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2026__A2
timestamp 1698431365
transform 1 0 20720 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2034__A2
timestamp 1698431365
transform -1 0 44464 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2036__S
timestamp 1698431365
transform 1 0 40432 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2037__B
timestamp 1698431365
transform 1 0 49056 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2051__A1
timestamp 1698431365
transform 1 0 48608 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2062__A1
timestamp 1698431365
transform 1 0 29792 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2062__B1
timestamp 1698431365
transform -1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2065__A1
timestamp 1698431365
transform -1 0 31808 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2067__A1
timestamp 1698431365
transform 1 0 27776 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2074__C
timestamp 1698431365
transform 1 0 31136 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2080__A1
timestamp 1698431365
transform -1 0 50624 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2080__B
timestamp 1698431365
transform 1 0 49952 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2096__A1
timestamp 1698431365
transform -1 0 50176 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2097__A1
timestamp 1698431365
transform 1 0 26992 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2099__A2
timestamp 1698431365
transform 1 0 28896 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2100__B2
timestamp 1698431365
transform 1 0 26208 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2101__A1
timestamp 1698431365
transform 1 0 30800 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2102__A3
timestamp 1698431365
transform 1 0 28560 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2108__A1
timestamp 1698431365
transform 1 0 31136 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2111__A2
timestamp 1698431365
transform 1 0 33152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2112__A1
timestamp 1698431365
transform 1 0 42672 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2117__A2
timestamp 1698431365
transform 1 0 34832 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2119__B
timestamp 1698431365
transform 1 0 24528 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2129__A1
timestamp 1698431365
transform 1 0 49840 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2132__A1
timestamp 1698431365
transform 1 0 24640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2134__B
timestamp 1698431365
transform -1 0 34384 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2137__A2
timestamp 1698431365
transform 1 0 28336 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2138__A2
timestamp 1698431365
transform 1 0 29904 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2139__A2
timestamp 1698431365
transform 1 0 30352 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2164__A2
timestamp 1698431365
transform 1 0 32480 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2171__I
timestamp 1698431365
transform 1 0 36736 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2187__A2
timestamp 1698431365
transform -1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2190__A1
timestamp 1698431365
transform -1 0 42448 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2190__C
timestamp 1698431365
transform 1 0 46704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2207__B2
timestamp 1698431365
transform 1 0 50288 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2216__B
timestamp 1698431365
transform 1 0 7168 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2223__I
timestamp 1698431365
transform -1 0 5712 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2228__A2
timestamp 1698431365
transform -1 0 6384 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2234__A1
timestamp 1698431365
transform -1 0 10640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2234__A2
timestamp 1698431365
transform 1 0 17472 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2234__C1
timestamp 1698431365
transform -1 0 9072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2238__I
timestamp 1698431365
transform 1 0 10080 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2244__B
timestamp 1698431365
transform -1 0 11312 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2249__C
timestamp 1698431365
transform 1 0 27776 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2255__A2
timestamp 1698431365
transform -1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2258__B
timestamp 1698431365
transform 1 0 16576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2261__A2
timestamp 1698431365
transform 1 0 30128 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2269__A1
timestamp 1698431365
transform 1 0 12208 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2269__B1
timestamp 1698431365
transform 1 0 12880 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2270__A1
timestamp 1698431365
transform 1 0 30576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2289__A2
timestamp 1698431365
transform -1 0 11424 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2289__B
timestamp 1698431365
transform -1 0 18256 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2291__I
timestamp 1698431365
transform 1 0 7504 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2292__I
timestamp 1698431365
transform 1 0 17472 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2294__A1
timestamp 1698431365
transform -1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2294__A3
timestamp 1698431365
transform -1 0 6720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2297__A1
timestamp 1698431365
transform 1 0 23744 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2297__A2
timestamp 1698431365
transform 1 0 25312 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2299__I
timestamp 1698431365
transform -1 0 5264 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2300__A2
timestamp 1698431365
transform -1 0 7056 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2300__A3
timestamp 1698431365
transform 1 0 12880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2303__A2
timestamp 1698431365
transform 1 0 9968 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2313__I
timestamp 1698431365
transform 1 0 44576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2322__A1
timestamp 1698431365
transform 1 0 16800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2322__A2
timestamp 1698431365
transform 1 0 15680 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2327__I0
timestamp 1698431365
transform 1 0 19376 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2327__I3
timestamp 1698431365
transform -1 0 19600 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2327__S1
timestamp 1698431365
transform 1 0 19824 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2330__A1
timestamp 1698431365
transform -1 0 10192 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2331__A1
timestamp 1698431365
transform 1 0 29232 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2331__A2
timestamp 1698431365
transform 1 0 27216 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2335__A2
timestamp 1698431365
transform -1 0 31248 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2339__A2
timestamp 1698431365
transform -1 0 15008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2339__B1
timestamp 1698431365
transform -1 0 16800 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2339__B2
timestamp 1698431365
transform -1 0 9072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2341__A1
timestamp 1698431365
transform 1 0 26768 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2343__A1
timestamp 1698431365
transform 1 0 21616 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2343__A2
timestamp 1698431365
transform 1 0 17584 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2350__A2
timestamp 1698431365
transform 1 0 27104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2359__A2
timestamp 1698431365
transform 1 0 8960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2362__A3
timestamp 1698431365
transform -1 0 8176 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2366__A1
timestamp 1698431365
transform 1 0 19824 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2367__A2
timestamp 1698431365
transform 1 0 5488 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2369__A2
timestamp 1698431365
transform 1 0 16800 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2370__A2
timestamp 1698431365
transform -1 0 6160 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2371__A3
timestamp 1698431365
transform -1 0 28448 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2373__A1
timestamp 1698431365
transform 1 0 25424 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2375__A2
timestamp 1698431365
transform -1 0 17696 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2378__A2
timestamp 1698431365
transform 1 0 13776 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2381__A2
timestamp 1698431365
transform 1 0 6944 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2382__A2
timestamp 1698431365
transform -1 0 21056 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2382__A3
timestamp 1698431365
transform -1 0 20272 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2384__I
timestamp 1698431365
transform 1 0 7280 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2385__A2
timestamp 1698431365
transform -1 0 17808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2387__I
timestamp 1698431365
transform -1 0 11424 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2391__C
timestamp 1698431365
transform -1 0 24528 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2392__A4
timestamp 1698431365
transform -1 0 31808 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2393__I
timestamp 1698431365
transform 1 0 38640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2395__A1
timestamp 1698431365
transform 1 0 9744 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2397__B
timestamp 1698431365
transform -1 0 15344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2398__A3
timestamp 1698431365
transform 1 0 27552 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2404__A2
timestamp 1698431365
transform -1 0 6496 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2405__A2
timestamp 1698431365
transform 1 0 13552 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2405__A3
timestamp 1698431365
transform 1 0 17472 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2407__A1
timestamp 1698431365
transform 1 0 4928 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2409__A1
timestamp 1698431365
transform -1 0 19936 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2413__B2
timestamp 1698431365
transform 1 0 31136 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2427__A1
timestamp 1698431365
transform -1 0 23072 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2430__A1
timestamp 1698431365
transform 1 0 20720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2430__A2
timestamp 1698431365
transform -1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2431__A1
timestamp 1698431365
transform 1 0 21392 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2436__I
timestamp 1698431365
transform 1 0 31472 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2437__A1
timestamp 1698431365
transform -1 0 7952 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2437__B
timestamp 1698431365
transform -1 0 10080 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2439__A2
timestamp 1698431365
transform 1 0 42336 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2444__A1
timestamp 1698431365
transform 1 0 13888 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2444__B1
timestamp 1698431365
transform 1 0 18592 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2444__B2
timestamp 1698431365
transform 1 0 15680 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2445__A1
timestamp 1698431365
transform 1 0 11872 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2445__A2
timestamp 1698431365
transform 1 0 12432 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2446__C
timestamp 1698431365
transform -1 0 13776 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2448__B
timestamp 1698431365
transform 1 0 16128 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2449__A3
timestamp 1698431365
transform 1 0 9744 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2450__A2
timestamp 1698431365
transform 1 0 12880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2451__A1
timestamp 1698431365
transform -1 0 20496 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2451__A2
timestamp 1698431365
transform 1 0 13552 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2453__A2
timestamp 1698431365
transform 1 0 38304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2454__A1
timestamp 1698431365
transform 1 0 20720 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2454__A2
timestamp 1698431365
transform 1 0 22960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2456__A2
timestamp 1698431365
transform -1 0 6720 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2457__A2
timestamp 1698431365
transform -1 0 8176 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2459__A1
timestamp 1698431365
transform 1 0 22400 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2459__B
timestamp 1698431365
transform 1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2460__A1
timestamp 1698431365
transform -1 0 8288 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2461__A1
timestamp 1698431365
transform -1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2461__A2
timestamp 1698431365
transform 1 0 27328 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2462__A3
timestamp 1698431365
transform -1 0 13328 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2463__A1
timestamp 1698431365
transform 1 0 29456 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2464__I
timestamp 1698431365
transform 1 0 31584 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2465__A2
timestamp 1698431365
transform -1 0 6608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2468__A2
timestamp 1698431365
transform 1 0 31136 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2473__A3
timestamp 1698431365
transform 1 0 32704 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2476__I0
timestamp 1698431365
transform -1 0 27776 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2476__S
timestamp 1698431365
transform 1 0 30352 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2477__A2
timestamp 1698431365
transform -1 0 30912 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2478__A1
timestamp 1698431365
transform 1 0 30240 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2487__A2
timestamp 1698431365
transform 1 0 38304 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2497__I
timestamp 1698431365
transform 1 0 25760 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2499__A2
timestamp 1698431365
transform -1 0 22624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2500__A1
timestamp 1698431365
transform 1 0 23520 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2501__I
timestamp 1698431365
transform -1 0 10976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2502__A1
timestamp 1698431365
transform -1 0 4816 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2502__B
timestamp 1698431365
transform -1 0 5600 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2503__A2
timestamp 1698431365
transform 1 0 9856 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2504__B1
timestamp 1698431365
transform -1 0 15904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2504__B2
timestamp 1698431365
transform 1 0 9856 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2507__A2
timestamp 1698431365
transform 1 0 16800 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2508__A1
timestamp 1698431365
transform 1 0 26320 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2508__B2
timestamp 1698431365
transform 1 0 21392 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2510__A2
timestamp 1698431365
transform 1 0 40992 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2511__A1
timestamp 1698431365
transform 1 0 42336 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2516__C
timestamp 1698431365
transform -1 0 6272 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2517__A1
timestamp 1698431365
transform -1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2518__A1
timestamp 1698431365
transform -1 0 6608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2518__A2
timestamp 1698431365
transform -1 0 6160 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2519__A1
timestamp 1698431365
transform -1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2520__A2
timestamp 1698431365
transform -1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2520__B
timestamp 1698431365
transform -1 0 6272 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2521__A1
timestamp 1698431365
transform -1 0 4368 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2525__A1
timestamp 1698431365
transform -1 0 8624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2525__B
timestamp 1698431365
transform -1 0 9520 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2526__A2
timestamp 1698431365
transform 1 0 6832 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2527__B
timestamp 1698431365
transform -1 0 7056 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2528__A1
timestamp 1698431365
transform -1 0 6048 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2529__A1
timestamp 1698431365
transform 1 0 31024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2530__A3
timestamp 1698431365
transform 1 0 31472 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2532__A3
timestamp 1698431365
transform 1 0 34272 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2533__A1
timestamp 1698431365
transform -1 0 30800 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2536__A2
timestamp 1698431365
transform -1 0 10192 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2537__A2
timestamp 1698431365
transform 1 0 19936 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2540__A3
timestamp 1698431365
transform 1 0 18368 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2547__A1
timestamp 1698431365
transform 1 0 46816 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2549__I
timestamp 1698431365
transform 1 0 43792 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2551__A1
timestamp 1698431365
transform 1 0 42336 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2561__A2
timestamp 1698431365
transform -1 0 11872 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2561__B
timestamp 1698431365
transform -1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2562__A1
timestamp 1698431365
transform -1 0 17696 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2562__A2
timestamp 1698431365
transform -1 0 18928 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2564__A2
timestamp 1698431365
transform 1 0 16240 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2565__A2
timestamp 1698431365
transform -1 0 18704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2566__A1
timestamp 1698431365
transform 1 0 15568 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2567__C
timestamp 1698431365
transform -1 0 21168 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2568__A1
timestamp 1698431365
transform -1 0 22624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2569__A2
timestamp 1698431365
transform 1 0 43008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2569__A3
timestamp 1698431365
transform 1 0 41552 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2571__A1
timestamp 1698431365
transform -1 0 41664 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2572__A1
timestamp 1698431365
transform -1 0 10528 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2575__B
timestamp 1698431365
transform -1 0 7168 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2575__C
timestamp 1698431365
transform -1 0 8736 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2576__A2
timestamp 1698431365
transform 1 0 24080 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2577__A1
timestamp 1698431365
transform 1 0 13664 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2585__A1
timestamp 1698431365
transform 1 0 43456 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2586__B
timestamp 1698431365
transform -1 0 10864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2588__A2
timestamp 1698431365
transform 1 0 28560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2588__B
timestamp 1698431365
transform 1 0 28112 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2589__A1
timestamp 1698431365
transform 1 0 26656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2589__A3
timestamp 1698431365
transform 1 0 27104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2597__I
timestamp 1698431365
transform 1 0 27664 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2598__I
timestamp 1698431365
transform 1 0 21840 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2600__A1
timestamp 1698431365
transform -1 0 9072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2600__B
timestamp 1698431365
transform -1 0 10080 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2601__I
timestamp 1698431365
transform -1 0 23520 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2602__A1
timestamp 1698431365
transform -1 0 25536 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2604__A2
timestamp 1698431365
transform -1 0 24416 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2609__A2
timestamp 1698431365
transform -1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2610__A2
timestamp 1698431365
transform -1 0 11984 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2611__A1
timestamp 1698431365
transform -1 0 12432 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2611__B2
timestamp 1698431365
transform -1 0 14448 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2631__A2
timestamp 1698431365
transform 1 0 14000 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2631__A3
timestamp 1698431365
transform 1 0 13104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2635__I
timestamp 1698431365
transform -1 0 23072 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2637__A2
timestamp 1698431365
transform 1 0 24304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2638__A1
timestamp 1698431365
transform -1 0 27328 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2638__A2
timestamp 1698431365
transform -1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2640__A1
timestamp 1698431365
transform 1 0 41664 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2642__A1
timestamp 1698431365
transform 1 0 44464 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2644__A1
timestamp 1698431365
transform 1 0 25088 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2644__A2
timestamp 1698431365
transform 1 0 25872 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2645__A2
timestamp 1698431365
transform 1 0 26320 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2646__A2
timestamp 1698431365
transform -1 0 20608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2649__A1
timestamp 1698431365
transform 1 0 23744 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2649__C
timestamp 1698431365
transform 1 0 26656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2667__B
timestamp 1698431365
transform 1 0 45024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2676__A1
timestamp 1698431365
transform 1 0 41664 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2680__A1
timestamp 1698431365
transform 1 0 22288 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2680__A2
timestamp 1698431365
transform 1 0 20720 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2680__C
timestamp 1698431365
transform -1 0 19040 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2682__I
timestamp 1698431365
transform 1 0 27328 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2689__I
timestamp 1698431365
transform -1 0 29568 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2691__A2
timestamp 1698431365
transform -1 0 21616 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2692__A1
timestamp 1698431365
transform 1 0 21280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2692__A2
timestamp 1698431365
transform -1 0 16576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2693__A2
timestamp 1698431365
transform -1 0 15344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2693__B2
timestamp 1698431365
transform -1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2694__A1
timestamp 1698431365
transform 1 0 14672 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2696__A1
timestamp 1698431365
transform 1 0 23072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2699__A2
timestamp 1698431365
transform -1 0 17360 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2699__A3
timestamp 1698431365
transform -1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2700__A2
timestamp 1698431365
transform -1 0 19824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2701__A1
timestamp 1698431365
transform -1 0 15456 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2702__A3
timestamp 1698431365
transform -1 0 22064 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2703__A2
timestamp 1698431365
transform 1 0 31584 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2706__A2
timestamp 1698431365
transform -1 0 38304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2722__A1
timestamp 1698431365
transform -1 0 11424 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2722__A2
timestamp 1698431365
transform 1 0 12656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2723__A2
timestamp 1698431365
transform -1 0 13776 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2724__A2
timestamp 1698431365
transform -1 0 15008 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2725__A3
timestamp 1698431365
transform -1 0 23968 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2731__A2
timestamp 1698431365
transform -1 0 14672 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2732__B
timestamp 1698431365
transform -1 0 5152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2733__B
timestamp 1698431365
transform -1 0 6720 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2734__B2
timestamp 1698431365
transform 1 0 22064 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2735__A2
timestamp 1698431365
transform 1 0 33824 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2736__A2
timestamp 1698431365
transform -1 0 33040 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2742__A2
timestamp 1698431365
transform 1 0 27552 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2744__A2
timestamp 1698431365
transform -1 0 18480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2745__A1
timestamp 1698431365
transform -1 0 19376 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2745__A2
timestamp 1698431365
transform -1 0 10976 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2746__A1
timestamp 1698431365
transform -1 0 24080 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2760__A2
timestamp 1698431365
transform -1 0 23968 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2760__A3
timestamp 1698431365
transform 1 0 27104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2762__B
timestamp 1698431365
transform -1 0 41216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2765__A1
timestamp 1698431365
transform -1 0 30688 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2767__A1
timestamp 1698431365
transform -1 0 26320 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2773__A1
timestamp 1698431365
transform 1 0 41216 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2776__S
timestamp 1698431365
transform 1 0 32368 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2788__A1
timestamp 1698431365
transform 1 0 29232 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2788__A2
timestamp 1698431365
transform 1 0 28560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2789__A1
timestamp 1698431365
transform 1 0 30240 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2789__A2
timestamp 1698431365
transform 1 0 31472 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2790__I0
timestamp 1698431365
transform -1 0 36848 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2791__I
timestamp 1698431365
transform -1 0 17696 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2792__A2
timestamp 1698431365
transform 1 0 19712 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2793__B
timestamp 1698431365
transform 1 0 20720 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2794__A1
timestamp 1698431365
transform 1 0 28784 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2794__A2
timestamp 1698431365
transform 1 0 29232 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2794__C
timestamp 1698431365
transform -1 0 28560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2798__A1
timestamp 1698431365
transform 1 0 28784 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2798__A2
timestamp 1698431365
transform 1 0 29232 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2798__B
timestamp 1698431365
transform 1 0 28224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2799__A1
timestamp 1698431365
transform 1 0 27776 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2803__C
timestamp 1698431365
transform 1 0 36064 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2817__A1
timestamp 1698431365
transform -1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2818__A2
timestamp 1698431365
transform 1 0 29232 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2822__A2
timestamp 1698431365
transform 1 0 35840 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2823__A1
timestamp 1698431365
transform 1 0 35168 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2823__C
timestamp 1698431365
transform 1 0 34720 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2837__A1
timestamp 1698431365
transform -1 0 22176 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2837__B
timestamp 1698431365
transform -1 0 23520 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2863__A1
timestamp 1698431365
transform 1 0 33936 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2864__I1
timestamp 1698431365
transform 1 0 33936 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2866__A1
timestamp 1698431365
transform 1 0 29680 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2867__I
timestamp 1698431365
transform 1 0 26208 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2871__A1
timestamp 1698431365
transform 1 0 9744 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2874__A2
timestamp 1698431365
transform -1 0 17696 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2875__A1
timestamp 1698431365
transform 1 0 18592 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2875__B1
timestamp 1698431365
transform 1 0 19264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2876__A2
timestamp 1698431365
transform -1 0 18704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2880__A1
timestamp 1698431365
transform -1 0 19264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2882__A1
timestamp 1698431365
transform 1 0 22288 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2883__A1
timestamp 1698431365
transform -1 0 20384 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2883__A2
timestamp 1698431365
transform 1 0 22736 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2884__A1
timestamp 1698431365
transform -1 0 22624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2885__A2
timestamp 1698431365
transform 1 0 22848 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2888__A2
timestamp 1698431365
transform 1 0 24192 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2888__B2
timestamp 1698431365
transform 1 0 24640 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2889__A1
timestamp 1698431365
transform 1 0 26208 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2892__A1
timestamp 1698431365
transform -1 0 22736 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2893__A1
timestamp 1698431365
transform 1 0 22960 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2894__A1
timestamp 1698431365
transform -1 0 18592 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2894__B1
timestamp 1698431365
transform -1 0 21616 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2895__A1
timestamp 1698431365
transform -1 0 20608 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2895__A2
timestamp 1698431365
transform -1 0 20832 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2897__A2
timestamp 1698431365
transform -1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2897__A3
timestamp 1698431365
transform 1 0 25872 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2900__A1
timestamp 1698431365
transform 1 0 23520 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2900__A2
timestamp 1698431365
transform -1 0 27664 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2902__A2
timestamp 1698431365
transform 1 0 23968 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2906__I1
timestamp 1698431365
transform -1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2908__A1
timestamp 1698431365
transform 1 0 43904 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2909__A1
timestamp 1698431365
transform 1 0 42336 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2913__CLK
timestamp 1698431365
transform 1 0 11760 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2914__CLK
timestamp 1698431365
transform 1 0 8848 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2915__CLK
timestamp 1698431365
transform 1 0 8736 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2916__CLK
timestamp 1698431365
transform -1 0 16688 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2919__CLK
timestamp 1698431365
transform 1 0 12544 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2920__CLK
timestamp 1698431365
transform 1 0 8288 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2921__CLK
timestamp 1698431365
transform 1 0 11312 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2922__CLK
timestamp 1698431365
transform 1 0 15232 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2923__CLK
timestamp 1698431365
transform 1 0 13552 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2929__D
timestamp 1698431365
transform 1 0 35728 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2929__RN
timestamp 1698431365
transform 1 0 30800 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2933__D
timestamp 1698431365
transform 1 0 40544 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2935__D
timestamp 1698431365
transform 1 0 43456 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_CLK_I
timestamp 1698431365
transform 1 0 18928 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout42_I
timestamp 1698431365
transform 1 0 40208 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout43_I
timestamp 1698431365
transform -1 0 39872 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout49_I
timestamp 1698431365
transform -1 0 35392 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout50_I
timestamp 1698431365
transform 1 0 14224 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout59_I
timestamp 1698431365
transform 1 0 10864 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout60_I
timestamp 1698431365
transform 1 0 30240 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout63_I
timestamp 1698431365
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout64_I
timestamp 1698431365
transform 1 0 43120 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout65_I
timestamp 1698431365
transform 1 0 28560 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 57680 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform 1 0 1792 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform 1 0 2464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output34_I
timestamp 1698431365
transform -1 0 4704 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output35_I
timestamp 1698431365
transform -1 0 28896 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output39_I
timestamp 1698431365
transform 1 0 4704 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output40_I
timestamp 1698431365
transform 1 0 4704 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output41_I
timestamp 1698431365
transform 1 0 36064 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19152 0 -1 31360
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_CLK
timestamp 1698431365
transform -1 0 17024 0 -1 32928
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_CLK
timestamp 1698431365
transform 1 0 26656 0 -1 31360
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout42
timestamp 1698431365
transform -1 0 39312 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout43
timestamp 1698431365
transform 1 0 38752 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout44
timestamp 1698431365
transform 1 0 39088 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout47
timestamp 1698431365
transform -1 0 39760 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout48
timestamp 1698431365
transform 1 0 39872 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout49
timestamp 1698431365
transform -1 0 31920 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout50
timestamp 1698431365
transform -1 0 15008 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout51
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout52
timestamp 1698431365
transform 1 0 11872 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout53
timestamp 1698431365
transform 1 0 15456 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout54
timestamp 1698431365
transform 1 0 7056 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout55
timestamp 1698431365
transform -1 0 10864 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout56
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout57
timestamp 1698431365
transform -1 0 8736 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout58
timestamp 1698431365
transform -1 0 9968 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout59
timestamp 1698431365
transform -1 0 10640 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout60
timestamp 1698431365
transform 1 0 29904 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout61
timestamp 1698431365
transform -1 0 43232 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout62
timestamp 1698431365
transform 1 0 43120 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout63
timestamp 1698431365
transform 1 0 37296 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout64
timestamp 1698431365
transform -1 0 44016 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout65
timestamp 1698431365
transform 1 0 29344 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout66
timestamp 1698431365
transform 1 0 7392 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_40 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5824 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_56 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7616 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_64 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8512 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_70 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_72 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_77
timestamp 1698431365
transform 1 0 9968 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_93
timestamp 1698431365
transform 1 0 11760 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_101
timestamp 1698431365
transform 1 0 12656 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_122
timestamp 1698431365
transform 1 0 15008 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_126
timestamp 1698431365
transform 1 0 15456 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_130
timestamp 1698431365
transform 1 0 15904 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_140
timestamp 1698431365
transform 1 0 17024 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_143
timestamp 1698431365
transform 1 0 17360 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_147
timestamp 1698431365
transform 1 0 17808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_151
timestamp 1698431365
transform 1 0 18256 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_155
timestamp 1698431365
transform 1 0 18704 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_161
timestamp 1698431365
transform 1 0 19376 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_165
timestamp 1698431365
transform 1 0 19824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_169
timestamp 1698431365
transform 1 0 20272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176
timestamp 1698431365
transform 1 0 21056 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_180
timestamp 1698431365
transform 1 0 21504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_182
timestamp 1698431365
transform 1 0 21728 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_185
timestamp 1698431365
transform 1 0 22064 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_189
timestamp 1698431365
transform 1 0 22512 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_191
timestamp 1698431365
transform 1 0 22736 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_194
timestamp 1698431365
transform 1 0 23072 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_198
timestamp 1698431365
transform 1 0 23520 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_202
timestamp 1698431365
transform 1 0 23968 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_287
timestamp 1698431365
transform 1 0 33488 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_303
timestamp 1698431365
transform 1 0 35280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_305
timestamp 1698431365
transform 1 0 35504 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_308
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_324
timestamp 1698431365
transform 1 0 37632 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_328
timestamp 1698431365
transform 1 0 38080 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_330
timestamp 1698431365
transform 1 0 38304 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_336
timestamp 1698431365
transform 1 0 38976 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_342
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_402
timestamp 1698431365
transform 1 0 46368 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_406
timestamp 1698431365
transform 1 0 46816 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_436
timestamp 1698431365
transform 1 0 50176 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_440
timestamp 1698431365
transform 1 0 50624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_474
timestamp 1698431365
transform 1 0 54432 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_478
timestamp 1698431365
transform 1 0 54880 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_494
timestamp 1698431365
transform 1 0 56672 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_502
timestamp 1698431365
transform 1 0 57568 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_506
timestamp 1698431365
transform 1 0 58016 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_508
timestamp 1698431365
transform 1 0 58240 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_104
timestamp 1698431365
transform 1 0 12992 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_112
timestamp 1698431365
transform 1 0 13888 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_114
timestamp 1698431365
transform 1 0 14112 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_117
timestamp 1698431365
transform 1 0 14448 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_121
timestamp 1698431365
transform 1 0 14896 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_125
timestamp 1698431365
transform 1 0 15344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_129
timestamp 1698431365
transform 1 0 15792 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_133
timestamp 1698431365
transform 1 0 16240 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_146
timestamp 1698431365
transform 1 0 17696 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_150
timestamp 1698431365
transform 1 0 18144 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_153
timestamp 1698431365
transform 1 0 18480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_168
timestamp 1698431365
transform 1 0 20160 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_172
timestamp 1698431365
transform 1 0 20608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_174
timestamp 1698431365
transform 1 0 20832 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_177
timestamp 1698431365
transform 1 0 21168 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_181
timestamp 1698431365
transform 1 0 21616 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_202
timestamp 1698431365
transform 1 0 23968 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_218
timestamp 1698431365
transform 1 0 25760 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_220
timestamp 1698431365
transform 1 0 25984 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_223
timestamp 1698431365
transform 1 0 26320 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_227
timestamp 1698431365
transform 1 0 26768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_229
timestamp 1698431365
transform 1 0 26992 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_232
timestamp 1698431365
transform 1 0 27328 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_240
timestamp 1698431365
transform 1 0 28224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_242
timestamp 1698431365
transform 1 0 28448 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_248
timestamp 1698431365
transform 1 0 29120 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_252
timestamp 1698431365
transform 1 0 29568 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_256
timestamp 1698431365
transform 1 0 30016 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698431365
transform 1 0 32480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_311
timestamp 1698431365
transform 1 0 36176 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_319
timestamp 1698431365
transform 1 0 37072 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_323
timestamp 1698431365
transform 1 0 37520 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_325
timestamp 1698431365
transform 1 0 37744 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_344
timestamp 1698431365
transform 1 0 39872 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_348
timestamp 1698431365
transform 1 0 40320 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_352
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_368
timestamp 1698431365
transform 1 0 42560 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_413
timestamp 1698431365
transform 1 0 47600 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_417
timestamp 1698431365
transform 1 0 48048 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_419
timestamp 1698431365
transform 1 0 48272 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_471
timestamp 1698431365
transform 1 0 54096 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_487
timestamp 1698431365
transform 1 0 55888 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_489
timestamp 1698431365
transform 1 0 56112 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_492
timestamp 1698431365
transform 1 0 56448 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_508
timestamp 1698431365
transform 1 0 58240 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_111
timestamp 1698431365
transform 1 0 13776 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_115
timestamp 1698431365
transform 1 0 14224 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_131
timestamp 1698431365
transform 1 0 16016 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_141
timestamp 1698431365
transform 1 0 17136 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_143
timestamp 1698431365
transform 1 0 17360 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_195
timestamp 1698431365
transform 1 0 23184 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_199
timestamp 1698431365
transform 1 0 23632 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_202
timestamp 1698431365
transform 1 0 23968 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_204
timestamp 1698431365
transform 1 0 24192 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_231
timestamp 1698431365
transform 1 0 27216 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_260
timestamp 1698431365
transform 1 0 30464 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_268
timestamp 1698431365
transform 1 0 31360 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_288
timestamp 1698431365
transform 1 0 33600 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_308
timestamp 1698431365
transform 1 0 35840 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_312
timestamp 1698431365
transform 1 0 36288 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_314
timestamp 1698431365
transform 1 0 36512 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_337
timestamp 1698431365
transform 1 0 39088 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_357
timestamp 1698431365
transform 1 0 41328 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_366
timestamp 1698431365
transform 1 0 42336 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_387
timestamp 1698431365
transform 1 0 44688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_413
timestamp 1698431365
transform 1 0 47600 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_436
timestamp 1698431365
transform 1 0 50176 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_448
timestamp 1698431365
transform 1 0 51520 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_452
timestamp 1698431365
transform 1 0 51968 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_454
timestamp 1698431365
transform 1 0 52192 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_457
timestamp 1698431365
transform 1 0 52528 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_489
timestamp 1698431365
transform 1 0 56112 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_505
timestamp 1698431365
transform 1 0 57904 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_88
timestamp 1698431365
transform 1 0 11200 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_92
timestamp 1698431365
transform 1 0 11648 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_95
timestamp 1698431365
transform 1 0 11984 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_99
timestamp 1698431365
transform 1 0 12432 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_103
timestamp 1698431365
transform 1 0 12880 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_113
timestamp 1698431365
transform 1 0 14000 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_144
timestamp 1698431365
transform 1 0 17472 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_183
timestamp 1698431365
transform 1 0 21840 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_187
timestamp 1698431365
transform 1 0 22288 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_201
timestamp 1698431365
transform 1 0 23856 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_203
timestamp 1698431365
transform 1 0 24080 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_206
timestamp 1698431365
transform 1 0 24416 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_220
timestamp 1698431365
transform 1 0 25984 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_222
timestamp 1698431365
transform 1 0 26208 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_258
timestamp 1698431365
transform 1 0 30240 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_262
timestamp 1698431365
transform 1 0 30688 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_266
timestamp 1698431365
transform 1 0 31136 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_273
timestamp 1698431365
transform 1 0 31920 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_277
timestamp 1698431365
transform 1 0 32368 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_279
timestamp 1698431365
transform 1 0 32592 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_298
timestamp 1698431365
transform 1 0 34720 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_302
timestamp 1698431365
transform 1 0 35168 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_326
timestamp 1698431365
transform 1 0 37856 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_347
timestamp 1698431365
transform 1 0 40208 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_349
timestamp 1698431365
transform 1 0 40432 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_368
timestamp 1698431365
transform 1 0 42560 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_389
timestamp 1698431365
transform 1 0 44912 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_394
timestamp 1698431365
transform 1 0 45472 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_398
timestamp 1698431365
transform 1 0 45920 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_445
timestamp 1698431365
transform 1 0 51184 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_477
timestamp 1698431365
transform 1 0 54768 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_485
timestamp 1698431365
transform 1 0 55664 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_489
timestamp 1698431365
transform 1 0 56112 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_492
timestamp 1698431365
transform 1 0 56448 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_508
timestamp 1698431365
transform 1 0 58240 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_69
timestamp 1698431365
transform 1 0 9072 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_73
timestamp 1698431365
transform 1 0 9520 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_75
timestamp 1698431365
transform 1 0 9744 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_78
timestamp 1698431365
transform 1 0 10080 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_86
timestamp 1698431365
transform 1 0 10976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_104
timestamp 1698431365
transform 1 0 12992 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_109
timestamp 1698431365
transform 1 0 13552 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_125
timestamp 1698431365
transform 1 0 15344 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_158
timestamp 1698431365
transform 1 0 19040 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_181
timestamp 1698431365
transform 1 0 21616 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_183
timestamp 1698431365
transform 1 0 21840 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_192
timestamp 1698431365
transform 1 0 22848 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_196
timestamp 1698431365
transform 1 0 23296 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_200
timestamp 1698431365
transform 1 0 23744 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_203
timestamp 1698431365
transform 1 0 24080 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_229
timestamp 1698431365
transform 1 0 26992 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_231
timestamp 1698431365
transform 1 0 27216 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_251
timestamp 1698431365
transform 1 0 29456 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_275
timestamp 1698431365
transform 1 0 32144 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_277
timestamp 1698431365
transform 1 0 32368 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698431365
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_323
timestamp 1698431365
transform 1 0 37520 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_340
timestamp 1698431365
transform 1 0 39424 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_372
timestamp 1698431365
transform 1 0 43008 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_380
timestamp 1698431365
transform 1 0 43904 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_384
timestamp 1698431365
transform 1 0 44352 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_387
timestamp 1698431365
transform 1 0 44688 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_403
timestamp 1698431365
transform 1 0 46480 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_411
timestamp 1698431365
transform 1 0 47376 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_429
timestamp 1698431365
transform 1 0 49392 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_445
timestamp 1698431365
transform 1 0 51184 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_453
timestamp 1698431365
transform 1 0 52080 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_457
timestamp 1698431365
transform 1 0 52528 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_489
timestamp 1698431365
transform 1 0 56112 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_505
timestamp 1698431365
transform 1 0 57904 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_170
timestamp 1698431365
transform 1 0 20384 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_186
timestamp 1698431365
transform 1 0 22176 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_190
timestamp 1698431365
transform 1 0 22624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_194
timestamp 1698431365
transform 1 0 23072 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_198
timestamp 1698431365
transform 1 0 23520 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_229
timestamp 1698431365
transform 1 0 26992 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_231
timestamp 1698431365
transform 1 0 27216 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_234
timestamp 1698431365
transform 1 0 27552 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_238
timestamp 1698431365
transform 1 0 28000 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_257
timestamp 1698431365
transform 1 0 30128 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_265
timestamp 1698431365
transform 1 0 31024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_284
timestamp 1698431365
transform 1 0 33152 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_308
timestamp 1698431365
transform 1 0 35840 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_312
timestamp 1698431365
transform 1 0 36288 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_344
timestamp 1698431365
transform 1 0 39872 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_348
timestamp 1698431365
transform 1 0 40320 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_352
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_383
timestamp 1698431365
transform 1 0 44240 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_391
timestamp 1698431365
transform 1 0 45136 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_410
timestamp 1698431365
transform 1 0 47264 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_418
timestamp 1698431365
transform 1 0 48160 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_422
timestamp 1698431365
transform 1 0 48608 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_434
timestamp 1698431365
transform 1 0 49952 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_448
timestamp 1698431365
transform 1 0 51520 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_480
timestamp 1698431365
transform 1 0 55104 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_488
timestamp 1698431365
transform 1 0 56000 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_492
timestamp 1698431365
transform 1 0 56448 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_500
timestamp 1698431365
transform 1 0 57344 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_504
timestamp 1698431365
transform 1 0 57792 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_69
timestamp 1698431365
transform 1 0 9072 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_77
timestamp 1698431365
transform 1 0 9968 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_81
timestamp 1698431365
transform 1 0 10416 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_83
timestamp 1698431365
transform 1 0 10640 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_86
timestamp 1698431365
transform 1 0 10976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_102
timestamp 1698431365
transform 1 0 12768 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_104
timestamp 1698431365
transform 1 0 12992 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_109
timestamp 1698431365
transform 1 0 13552 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_128
timestamp 1698431365
transform 1 0 15680 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_134
timestamp 1698431365
transform 1 0 16352 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_181
timestamp 1698431365
transform 1 0 21616 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_183
timestamp 1698431365
transform 1 0 21840 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_217
timestamp 1698431365
transform 1 0 25648 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_221
timestamp 1698431365
transform 1 0 26096 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_225
timestamp 1698431365
transform 1 0 26544 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_260
timestamp 1698431365
transform 1 0 30464 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_268
timestamp 1698431365
transform 1 0 31360 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_272
timestamp 1698431365
transform 1 0 31808 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_287
timestamp 1698431365
transform 1 0 33488 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_295
timestamp 1698431365
transform 1 0 34384 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_299
timestamp 1698431365
transform 1 0 34832 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_312
timestamp 1698431365
transform 1 0 36288 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_314
timestamp 1698431365
transform 1 0 36512 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_325
timestamp 1698431365
transform 1 0 37744 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_329
timestamp 1698431365
transform 1 0 38192 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_331
timestamp 1698431365
transform 1 0 38416 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_337
timestamp 1698431365
transform 1 0 39088 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_353
timestamp 1698431365
transform 1 0 40880 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_375
timestamp 1698431365
transform 1 0 43344 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_383
timestamp 1698431365
transform 1 0 44240 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_401
timestamp 1698431365
transform 1 0 46256 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_454
timestamp 1698431365
transform 1 0 52192 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_457
timestamp 1698431365
transform 1 0 52528 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_473
timestamp 1698431365
transform 1 0 54320 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_481
timestamp 1698431365
transform 1 0 55216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698431365
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_78
timestamp 1698431365
transform 1 0 10080 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_82
timestamp 1698431365
transform 1 0 10528 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_86
timestamp 1698431365
transform 1 0 10976 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_90
timestamp 1698431365
transform 1 0 11424 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_103
timestamp 1698431365
transform 1 0 12880 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_105
timestamp 1698431365
transform 1 0 13104 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_118
timestamp 1698431365
transform 1 0 14560 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_199
timestamp 1698431365
transform 1 0 23632 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_228
timestamp 1698431365
transform 1 0 26880 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_232
timestamp 1698431365
transform 1 0 27328 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_242
timestamp 1698431365
transform 1 0 28448 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_244
timestamp 1698431365
transform 1 0 28672 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_247
timestamp 1698431365
transform 1 0 29008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_251
timestamp 1698431365
transform 1 0 29456 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_255
timestamp 1698431365
transform 1 0 29904 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_263
timestamp 1698431365
transform 1 0 30800 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_267
timestamp 1698431365
transform 1 0 31248 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_313
timestamp 1698431365
transform 1 0 36400 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_317
timestamp 1698431365
transform 1 0 36848 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_325
timestamp 1698431365
transform 1 0 37744 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_327
timestamp 1698431365
transform 1 0 37968 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698431365
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_352
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_356
timestamp 1698431365
transform 1 0 41216 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_358
timestamp 1698431365
transform 1 0 41440 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_375
timestamp 1698431365
transform 1 0 43344 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_383
timestamp 1698431365
transform 1 0 44240 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_402
timestamp 1698431365
transform 1 0 46368 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_418
timestamp 1698431365
transform 1 0 48160 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_422
timestamp 1698431365
transform 1 0 48608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_424
timestamp 1698431365
transform 1 0 48832 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_450
timestamp 1698431365
transform 1 0 51744 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_482
timestamp 1698431365
transform 1 0 55328 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_492
timestamp 1698431365
transform 1 0 56448 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_508
timestamp 1698431365
transform 1 0 58240 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_53
timestamp 1698431365
transform 1 0 7280 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_61
timestamp 1698431365
transform 1 0 8176 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_65
timestamp 1698431365
transform 1 0 8624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_69
timestamp 1698431365
transform 1 0 9072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_100
timestamp 1698431365
transform 1 0 12544 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_102
timestamp 1698431365
transform 1 0 12768 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_131
timestamp 1698431365
transform 1 0 16016 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_147
timestamp 1698431365
transform 1 0 17808 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_165
timestamp 1698431365
transform 1 0 19824 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_193
timestamp 1698431365
transform 1 0 22960 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_207
timestamp 1698431365
transform 1 0 24528 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_211
timestamp 1698431365
transform 1 0 24976 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_226
timestamp 1698431365
transform 1 0 26656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_237
timestamp 1698431365
transform 1 0 27888 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_243
timestamp 1698431365
transform 1 0 28560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_255
timestamp 1698431365
transform 1 0 29904 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_271
timestamp 1698431365
transform 1 0 31696 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_275
timestamp 1698431365
transform 1 0 32144 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_279
timestamp 1698431365
transform 1 0 32592 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_283
timestamp 1698431365
transform 1 0 33040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_299
timestamp 1698431365
transform 1 0 34832 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_303
timestamp 1698431365
transform 1 0 35280 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_305
timestamp 1698431365
transform 1 0 35504 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_310
timestamp 1698431365
transform 1 0 36064 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_314
timestamp 1698431365
transform 1 0 36512 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_325
timestamp 1698431365
transform 1 0 37744 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_327
timestamp 1698431365
transform 1 0 37968 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_359
timestamp 1698431365
transform 1 0 41552 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_375
timestamp 1698431365
transform 1 0 43344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_387
timestamp 1698431365
transform 1 0 44688 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_417
timestamp 1698431365
transform 1 0 48048 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_421
timestamp 1698431365
transform 1 0 48496 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_423
timestamp 1698431365
transform 1 0 48720 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_430
timestamp 1698431365
transform 1 0 49504 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_446
timestamp 1698431365
transform 1 0 51296 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_454
timestamp 1698431365
transform 1 0 52192 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_457
timestamp 1698431365
transform 1 0 52528 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_489
timestamp 1698431365
transform 1 0 56112 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_34
timestamp 1698431365
transform 1 0 5152 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_50
timestamp 1698431365
transform 1 0 6944 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_58
timestamp 1698431365
transform 1 0 7840 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_62
timestamp 1698431365
transform 1 0 8288 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_66
timestamp 1698431365
transform 1 0 8736 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_74
timestamp 1698431365
transform 1 0 9632 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_120
timestamp 1698431365
transform 1 0 14784 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_135
timestamp 1698431365
transform 1 0 16464 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_137
timestamp 1698431365
transform 1 0 16688 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_164
timestamp 1698431365
transform 1 0 19712 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_191
timestamp 1698431365
transform 1 0 22736 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_195
timestamp 1698431365
transform 1 0 23184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_197
timestamp 1698431365
transform 1 0 23408 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_207
timestamp 1698431365
transform 1 0 24528 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_209
timestamp 1698431365
transform 1 0 24752 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_216
timestamp 1698431365
transform 1 0 25536 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_220
timestamp 1698431365
transform 1 0 25984 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_222
timestamp 1698431365
transform 1 0 26208 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_240
timestamp 1698431365
transform 1 0 28224 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_244
timestamp 1698431365
transform 1 0 28672 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_247
timestamp 1698431365
transform 1 0 29008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_251
timestamp 1698431365
transform 1 0 29456 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_253
timestamp 1698431365
transform 1 0 29680 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_277
timestamp 1698431365
transform 1 0 32368 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_279
timestamp 1698431365
transform 1 0 32592 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_305
timestamp 1698431365
transform 1 0 35504 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_307
timestamp 1698431365
transform 1 0 35728 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_313
timestamp 1698431365
transform 1 0 36400 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_317
timestamp 1698431365
transform 1 0 36848 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_319
timestamp 1698431365
transform 1 0 37072 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_328
timestamp 1698431365
transform 1 0 38080 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_342
timestamp 1698431365
transform 1 0 39648 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_358
timestamp 1698431365
transform 1 0 41440 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_374
timestamp 1698431365
transform 1 0 43232 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_390
timestamp 1698431365
transform 1 0 45024 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_398
timestamp 1698431365
transform 1 0 45920 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_415
timestamp 1698431365
transform 1 0 47824 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_419
timestamp 1698431365
transform 1 0 48272 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_439
timestamp 1698431365
transform 1 0 50512 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_471
timestamp 1698431365
transform 1 0 54096 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_487
timestamp 1698431365
transform 1 0 55888 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_489
timestamp 1698431365
transform 1 0 56112 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_492
timestamp 1698431365
transform 1 0 56448 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_500
timestamp 1698431365
transform 1 0 57344 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_53
timestamp 1698431365
transform 1 0 7280 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_57
timestamp 1698431365
transform 1 0 7728 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_77
timestamp 1698431365
transform 1 0 9968 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_96
timestamp 1698431365
transform 1 0 12096 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_169
timestamp 1698431365
transform 1 0 20272 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_179
timestamp 1698431365
transform 1 0 21392 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_196
timestamp 1698431365
transform 1 0 23296 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_220
timestamp 1698431365
transform 1 0 25984 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_222
timestamp 1698431365
transform 1 0 26208 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_239
timestamp 1698431365
transform 1 0 28112 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_270
timestamp 1698431365
transform 1 0 31584 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_278
timestamp 1698431365
transform 1 0 32480 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_280
timestamp 1698431365
transform 1 0 32704 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_306
timestamp 1698431365
transform 1 0 35616 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_314
timestamp 1698431365
transform 1 0 36512 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_330
timestamp 1698431365
transform 1 0 38304 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_338
timestamp 1698431365
transform 1 0 39200 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_352
timestamp 1698431365
transform 1 0 40768 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_356
timestamp 1698431365
transform 1 0 41216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_363
timestamp 1698431365
transform 1 0 42000 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_383
timestamp 1698431365
transform 1 0 44240 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_387
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_399
timestamp 1698431365
transform 1 0 46032 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_417
timestamp 1698431365
transform 1 0 48048 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_451
timestamp 1698431365
transform 1 0 51856 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_457
timestamp 1698431365
transform 1 0 52528 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_473
timestamp 1698431365
transform 1 0 54320 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_481
timestamp 1698431365
transform 1 0 55216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_34
timestamp 1698431365
transform 1 0 5152 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_42
timestamp 1698431365
transform 1 0 6048 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_48
timestamp 1698431365
transform 1 0 6720 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_68
timestamp 1698431365
transform 1 0 8960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_103
timestamp 1698431365
transform 1 0 12880 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_133
timestamp 1698431365
transform 1 0 16240 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_137
timestamp 1698431365
transform 1 0 16688 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_186
timestamp 1698431365
transform 1 0 22176 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_196
timestamp 1698431365
transform 1 0 23296 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_208
timestamp 1698431365
transform 1 0 24640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_216
timestamp 1698431365
transform 1 0 25536 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_218
timestamp 1698431365
transform 1 0 25760 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_224
timestamp 1698431365
transform 1 0 26432 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_228
timestamp 1698431365
transform 1 0 26880 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_247
timestamp 1698431365
transform 1 0 29008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_256
timestamp 1698431365
transform 1 0 30016 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_267
timestamp 1698431365
transform 1 0 31248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_271
timestamp 1698431365
transform 1 0 31696 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_279
timestamp 1698431365
transform 1 0 32592 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_288
timestamp 1698431365
transform 1 0 33600 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_292
timestamp 1698431365
transform 1 0 34048 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_296
timestamp 1698431365
transform 1 0 34496 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_300
timestamp 1698431365
transform 1 0 34944 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_304
timestamp 1698431365
transform 1 0 35392 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_324
timestamp 1698431365
transform 1 0 37632 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_328
timestamp 1698431365
transform 1 0 38080 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_344
timestamp 1698431365
transform 1 0 39872 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_348
timestamp 1698431365
transform 1 0 40320 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_352
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_370
timestamp 1698431365
transform 1 0 42784 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_383
timestamp 1698431365
transform 1 0 44240 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_387
timestamp 1698431365
transform 1 0 44688 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_395
timestamp 1698431365
transform 1 0 45584 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_399
timestamp 1698431365
transform 1 0 46032 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_414
timestamp 1698431365
transform 1 0 47712 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_418
timestamp 1698431365
transform 1 0 48160 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_422
timestamp 1698431365
transform 1 0 48608 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_430
timestamp 1698431365
transform 1 0 49504 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_442
timestamp 1698431365
transform 1 0 50848 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_474
timestamp 1698431365
transform 1 0 54432 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_492
timestamp 1698431365
transform 1 0 56448 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_508
timestamp 1698431365
transform 1 0 58240 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_47
timestamp 1698431365
transform 1 0 6608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_51
timestamp 1698431365
transform 1 0 7056 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_55
timestamp 1698431365
transform 1 0 7504 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_101
timestamp 1698431365
transform 1 0 12656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_109
timestamp 1698431365
transform 1 0 13552 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_139
timestamp 1698431365
transform 1 0 16912 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_173
timestamp 1698431365
transform 1 0 20720 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_179
timestamp 1698431365
transform 1 0 21392 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_241
timestamp 1698431365
transform 1 0 28336 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_262
timestamp 1698431365
transform 1 0 30688 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_264
timestamp 1698431365
transform 1 0 30912 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_267
timestamp 1698431365
transform 1 0 31248 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_271
timestamp 1698431365
transform 1 0 31696 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_273
timestamp 1698431365
transform 1 0 31920 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_280
timestamp 1698431365
transform 1 0 32704 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_296
timestamp 1698431365
transform 1 0 34496 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_304
timestamp 1698431365
transform 1 0 35392 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_349
timestamp 1698431365
transform 1 0 40432 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_357
timestamp 1698431365
transform 1 0 41328 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_378
timestamp 1698431365
transform 1 0 43680 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_382
timestamp 1698431365
transform 1 0 44128 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_384
timestamp 1698431365
transform 1 0 44352 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_387
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_419
timestamp 1698431365
transform 1 0 48272 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_423
timestamp 1698431365
transform 1 0 48720 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_445
timestamp 1698431365
transform 1 0 51184 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_453
timestamp 1698431365
transform 1 0 52080 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_457
timestamp 1698431365
transform 1 0 52528 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_489
timestamp 1698431365
transform 1 0 56112 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_34
timestamp 1698431365
transform 1 0 5152 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_44
timestamp 1698431365
transform 1 0 6272 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_64
timestamp 1698431365
transform 1 0 8512 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_134
timestamp 1698431365
transform 1 0 16352 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_197
timestamp 1698431365
transform 1 0 23408 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_208
timestamp 1698431365
transform 1 0 24640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_222
timestamp 1698431365
transform 1 0 26208 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_275
timestamp 1698431365
transform 1 0 32144 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_279
timestamp 1698431365
transform 1 0 32592 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_305
timestamp 1698431365
transform 1 0 35504 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_313
timestamp 1698431365
transform 1 0 36400 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_342
timestamp 1698431365
transform 1 0 39648 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_368
timestamp 1698431365
transform 1 0 42560 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_372
timestamp 1698431365
transform 1 0 43008 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_379
timestamp 1698431365
transform 1 0 43792 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_414
timestamp 1698431365
transform 1 0 47712 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_418
timestamp 1698431365
transform 1 0 48160 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_422
timestamp 1698431365
transform 1 0 48608 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_461
timestamp 1698431365
transform 1 0 52976 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_477
timestamp 1698431365
transform 1 0 54768 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_485
timestamp 1698431365
transform 1 0 55664 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_489
timestamp 1698431365
transform 1 0 56112 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_492
timestamp 1698431365
transform 1 0 56448 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_500
timestamp 1698431365
transform 1 0 57344 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_504
timestamp 1698431365
transform 1 0 57792 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_18
timestamp 1698431365
transform 1 0 3360 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_26
timestamp 1698431365
transform 1 0 4256 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_30
timestamp 1698431365
transform 1 0 4704 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_32
timestamp 1698431365
transform 1 0 4928 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_41
timestamp 1698431365
transform 1 0 5936 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_44
timestamp 1698431365
transform 1 0 6272 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_203
timestamp 1698431365
transform 1 0 24080 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_253
timestamp 1698431365
transform 1 0 29680 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_286
timestamp 1698431365
transform 1 0 33376 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_314
timestamp 1698431365
transform 1 0 36512 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_321
timestamp 1698431365
transform 1 0 37296 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_323
timestamp 1698431365
transform 1 0 37520 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_350
timestamp 1698431365
transform 1 0 40544 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_354
timestamp 1698431365
transform 1 0 40992 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_403
timestamp 1698431365
transform 1 0 46480 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_405
timestamp 1698431365
transform 1 0 46704 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_435
timestamp 1698431365
transform 1 0 50064 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_451
timestamp 1698431365
transform 1 0 51856 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_457
timestamp 1698431365
transform 1 0 52528 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_473
timestamp 1698431365
transform 1 0 54320 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_481
timestamp 1698431365
transform 1 0 55216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_18
timestamp 1698431365
transform 1 0 3360 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_26
timestamp 1698431365
transform 1 0 4256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_30
timestamp 1698431365
transform 1 0 4704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_34
timestamp 1698431365
transform 1 0 5152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_38
timestamp 1698431365
transform 1 0 5600 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_42
timestamp 1698431365
transform 1 0 6048 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_80
timestamp 1698431365
transform 1 0 10304 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_82
timestamp 1698431365
transform 1 0 10528 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_85
timestamp 1698431365
transform 1 0 10864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_161
timestamp 1698431365
transform 1 0 19376 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_231
timestamp 1698431365
transform 1 0 27216 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_233
timestamp 1698431365
transform 1 0 27440 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_259
timestamp 1698431365
transform 1 0 30352 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_273
timestamp 1698431365
transform 1 0 31920 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_277
timestamp 1698431365
transform 1 0 32368 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698431365
transform 1 0 32592 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_305
timestamp 1698431365
transform 1 0 35504 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_313
timestamp 1698431365
transform 1 0 36400 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_317
timestamp 1698431365
transform 1 0 36848 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_357
timestamp 1698431365
transform 1 0 41328 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_361
timestamp 1698431365
transform 1 0 41776 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_370
timestamp 1698431365
transform 1 0 42784 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_374
timestamp 1698431365
transform 1 0 43232 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_378
timestamp 1698431365
transform 1 0 43680 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_386
timestamp 1698431365
transform 1 0 44576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_399
timestamp 1698431365
transform 1 0 46032 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_422
timestamp 1698431365
transform 1 0 48608 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_438
timestamp 1698431365
transform 1 0 50400 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_466
timestamp 1698431365
transform 1 0 53536 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_482
timestamp 1698431365
transform 1 0 55328 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_492
timestamp 1698431365
transform 1 0 56448 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_508
timestamp 1698431365
transform 1 0 58240 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_18
timestamp 1698431365
transform 1 0 3360 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_22
timestamp 1698431365
transform 1 0 3808 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_24
timestamp 1698431365
transform 1 0 4032 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_27
timestamp 1698431365
transform 1 0 4368 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_31
timestamp 1698431365
transform 1 0 4816 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_62
timestamp 1698431365
transform 1 0 8288 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_133
timestamp 1698431365
transform 1 0 16240 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_173
timestamp 1698431365
transform 1 0 20720 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_242
timestamp 1698431365
transform 1 0 28448 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698431365
transform 1 0 28672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_256
timestamp 1698431365
transform 1 0 30016 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_260
timestamp 1698431365
transform 1 0 30464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_264
timestamp 1698431365
transform 1 0 30912 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_268
timestamp 1698431365
transform 1 0 31360 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_272
timestamp 1698431365
transform 1 0 31808 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_280
timestamp 1698431365
transform 1 0 32704 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_290
timestamp 1698431365
transform 1 0 33824 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_292
timestamp 1698431365
transform 1 0 34048 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_312
timestamp 1698431365
transform 1 0 36288 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_314
timestamp 1698431365
transform 1 0 36512 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_340
timestamp 1698431365
transform 1 0 39424 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_364
timestamp 1698431365
transform 1 0 42112 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_368
timestamp 1698431365
transform 1 0 42560 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_384
timestamp 1698431365
transform 1 0 44352 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_387
timestamp 1698431365
transform 1 0 44688 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_419
timestamp 1698431365
transform 1 0 48272 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_427
timestamp 1698431365
transform 1 0 49168 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_431
timestamp 1698431365
transform 1 0 49616 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_450
timestamp 1698431365
transform 1 0 51744 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_454
timestamp 1698431365
transform 1 0 52192 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_463
timestamp 1698431365
transform 1 0 53200 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_479
timestamp 1698431365
transform 1 0 54992 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_18
timestamp 1698431365
transform 1 0 3360 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_26
timestamp 1698431365
transform 1 0 4256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_30
timestamp 1698431365
transform 1 0 4704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_32
timestamp 1698431365
transform 1 0 4928 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_35
timestamp 1698431365
transform 1 0 5264 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_39
timestamp 1698431365
transform 1 0 5712 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_43
timestamp 1698431365
transform 1 0 6160 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_47
timestamp 1698431365
transform 1 0 6608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_67
timestamp 1698431365
transform 1 0 8848 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_69
timestamp 1698431365
transform 1 0 9072 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_76
timestamp 1698431365
transform 1 0 9856 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_79
timestamp 1698431365
transform 1 0 10192 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_239
timestamp 1698431365
transform 1 0 28112 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_286
timestamp 1698431365
transform 1 0 33376 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_288
timestamp 1698431365
transform 1 0 33600 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_329
timestamp 1698431365
transform 1 0 38192 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_345
timestamp 1698431365
transform 1 0 39984 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_349
timestamp 1698431365
transform 1 0 40432 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_377
timestamp 1698431365
transform 1 0 43568 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_381
timestamp 1698431365
transform 1 0 44016 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_389
timestamp 1698431365
transform 1 0 44912 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_391
timestamp 1698431365
transform 1 0 45136 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_411
timestamp 1698431365
transform 1 0 47376 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_419
timestamp 1698431365
transform 1 0 48272 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_422
timestamp 1698431365
transform 1 0 48608 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_430
timestamp 1698431365
transform 1 0 49504 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_432
timestamp 1698431365
transform 1 0 49728 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_469
timestamp 1698431365
transform 1 0 53872 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_485
timestamp 1698431365
transform 1 0 55664 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_489
timestamp 1698431365
transform 1 0 56112 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_492
timestamp 1698431365
transform 1 0 56448 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_500
timestamp 1698431365
transform 1 0 57344 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_504
timestamp 1698431365
transform 1 0 57792 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_6
timestamp 1698431365
transform 1 0 2016 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_14
timestamp 1698431365
transform 1 0 2912 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_18
timestamp 1698431365
transform 1 0 3360 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_20
timestamp 1698431365
transform 1 0 3584 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_104
timestamp 1698431365
transform 1 0 12992 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_182
timestamp 1698431365
transform 1 0 21728 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_197
timestamp 1698431365
transform 1 0 23408 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_199
timestamp 1698431365
transform 1 0 23632 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_249
timestamp 1698431365
transform 1 0 29232 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_288
timestamp 1698431365
transform 1 0 33600 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_292
timestamp 1698431365
transform 1 0 34048 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_312
timestamp 1698431365
transform 1 0 36288 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_314
timestamp 1698431365
transform 1 0 36512 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_339
timestamp 1698431365
transform 1 0 39312 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_355
timestamp 1698431365
transform 1 0 41104 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_367
timestamp 1698431365
transform 1 0 42448 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_382
timestamp 1698431365
transform 1 0 44128 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_384
timestamp 1698431365
transform 1 0 44352 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_387
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_391
timestamp 1698431365
transform 1 0 45136 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_451
timestamp 1698431365
transform 1 0 51856 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_457
timestamp 1698431365
transform 1 0 52528 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_473
timestamp 1698431365
transform 1 0 54320 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_481
timestamp 1698431365
transform 1 0 55216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_18
timestamp 1698431365
transform 1 0 3360 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_26
timestamp 1698431365
transform 1 0 4256 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_30
timestamp 1698431365
transform 1 0 4704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_36
timestamp 1698431365
transform 1 0 5376 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_40
timestamp 1698431365
transform 1 0 5824 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_43
timestamp 1698431365
transform 1 0 6160 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_47
timestamp 1698431365
transform 1 0 6608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_69
timestamp 1698431365
transform 1 0 9072 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_74
timestamp 1698431365
transform 1 0 9632 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_121
timestamp 1698431365
transform 1 0 14896 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_138
timestamp 1698431365
transform 1 0 16800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_148
timestamp 1698431365
transform 1 0 17920 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_185
timestamp 1698431365
transform 1 0 22064 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_187
timestamp 1698431365
transform 1 0 22288 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_205
timestamp 1698431365
transform 1 0 24304 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_207
timestamp 1698431365
transform 1 0 24528 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_222
timestamp 1698431365
transform 1 0 26208 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_228
timestamp 1698431365
transform 1 0 26880 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_232
timestamp 1698431365
transform 1 0 27328 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_244
timestamp 1698431365
transform 1 0 28672 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_246
timestamp 1698431365
transform 1 0 28896 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_272
timestamp 1698431365
transform 1 0 31808 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_298
timestamp 1698431365
transform 1 0 34720 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_300
timestamp 1698431365
transform 1 0 34944 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_327
timestamp 1698431365
transform 1 0 37968 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_329
timestamp 1698431365
transform 1 0 38192 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_348
timestamp 1698431365
transform 1 0 40320 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_352
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_368
timestamp 1698431365
transform 1 0 42560 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_372
timestamp 1698431365
transform 1 0 43008 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_383
timestamp 1698431365
transform 1 0 44240 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_391
timestamp 1698431365
transform 1 0 45136 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_395
timestamp 1698431365
transform 1 0 45584 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_404
timestamp 1698431365
transform 1 0 46592 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_408
timestamp 1698431365
transform 1 0 47040 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_414
timestamp 1698431365
transform 1 0 47712 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_418
timestamp 1698431365
transform 1 0 48160 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_422
timestamp 1698431365
transform 1 0 48608 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_443
timestamp 1698431365
transform 1 0 50960 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_475
timestamp 1698431365
transform 1 0 54544 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_483
timestamp 1698431365
transform 1 0 55440 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_487
timestamp 1698431365
transform 1 0 55888 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_489
timestamp 1698431365
transform 1 0 56112 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_492
timestamp 1698431365
transform 1 0 56448 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_508
timestamp 1698431365
transform 1 0 58240 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_43
timestamp 1698431365
transform 1 0 6160 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_63
timestamp 1698431365
transform 1 0 8400 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_77
timestamp 1698431365
transform 1 0 9968 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_150
timestamp 1698431365
transform 1 0 18144 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_173
timestamp 1698431365
transform 1 0 20720 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_207
timestamp 1698431365
transform 1 0 24528 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_209
timestamp 1698431365
transform 1 0 24752 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_228
timestamp 1698431365
transform 1 0 26880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_232
timestamp 1698431365
transform 1 0 27328 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_236
timestamp 1698431365
transform 1 0 27776 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_238
timestamp 1698431365
transform 1 0 28000 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_241
timestamp 1698431365
transform 1 0 28336 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_257
timestamp 1698431365
transform 1 0 30128 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_261
timestamp 1698431365
transform 1 0 30576 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_265
timestamp 1698431365
transform 1 0 31024 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_268
timestamp 1698431365
transform 1 0 31360 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_272
timestamp 1698431365
transform 1 0 31808 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_282
timestamp 1698431365
transform 1 0 32928 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_286
timestamp 1698431365
transform 1 0 33376 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_293
timestamp 1698431365
transform 1 0 34160 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_301
timestamp 1698431365
transform 1 0 35056 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_305
timestamp 1698431365
transform 1 0 35504 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_337
timestamp 1698431365
transform 1 0 39088 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_341
timestamp 1698431365
transform 1 0 39536 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_353
timestamp 1698431365
transform 1 0 40880 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_361
timestamp 1698431365
transform 1 0 41776 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_365
timestamp 1698431365
transform 1 0 42224 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_368
timestamp 1698431365
transform 1 0 42560 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_372
timestamp 1698431365
transform 1 0 43008 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_387
timestamp 1698431365
transform 1 0 44688 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_395
timestamp 1698431365
transform 1 0 45584 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_399
timestamp 1698431365
transform 1 0 46032 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_408
timestamp 1698431365
transform 1 0 47040 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_463
timestamp 1698431365
transform 1 0 53200 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_495
timestamp 1698431365
transform 1 0 56784 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_503
timestamp 1698431365
transform 1 0 57680 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_18
timestamp 1698431365
transform 1 0 3360 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_26
timestamp 1698431365
transform 1 0 4256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_30
timestamp 1698431365
transform 1 0 4704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_42
timestamp 1698431365
transform 1 0 6048 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_81
timestamp 1698431365
transform 1 0 10416 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_138
timestamp 1698431365
transform 1 0 16800 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_151
timestamp 1698431365
transform 1 0 18256 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_199
timestamp 1698431365
transform 1 0 23632 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_201
timestamp 1698431365
transform 1 0 23856 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_229
timestamp 1698431365
transform 1 0 26992 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_265
timestamp 1698431365
transform 1 0 31024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_267
timestamp 1698431365
transform 1 0 31248 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_277
timestamp 1698431365
transform 1 0 32368 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698431365
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_301
timestamp 1698431365
transform 1 0 35056 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_305
timestamp 1698431365
transform 1 0 35504 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_321
timestamp 1698431365
transform 1 0 37296 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_325
timestamp 1698431365
transform 1 0 37744 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_334
timestamp 1698431365
transform 1 0 38752 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_336
timestamp 1698431365
transform 1 0 38976 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_352
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_422
timestamp 1698431365
transform 1 0 48608 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_431
timestamp 1698431365
transform 1 0 49616 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_463
timestamp 1698431365
transform 1 0 53200 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_479
timestamp 1698431365
transform 1 0 54992 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_487
timestamp 1698431365
transform 1 0 55888 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_489
timestamp 1698431365
transform 1 0 56112 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_492
timestamp 1698431365
transform 1 0 56448 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_500
timestamp 1698431365
transform 1 0 57344 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_504
timestamp 1698431365
transform 1 0 57792 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_41
timestamp 1698431365
transform 1 0 5936 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_75
timestamp 1698431365
transform 1 0 9744 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_77
timestamp 1698431365
transform 1 0 9968 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_152
timestamp 1698431365
transform 1 0 18368 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_156
timestamp 1698431365
transform 1 0 18816 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_158
timestamp 1698431365
transform 1 0 19040 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_249
timestamp 1698431365
transform 1 0 29232 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_283
timestamp 1698431365
transform 1 0 33040 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_285
timestamp 1698431365
transform 1 0 33264 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698431365
transform 1 0 37296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_331
timestamp 1698431365
transform 1 0 38416 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_335
timestamp 1698431365
transform 1 0 38864 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_339
timestamp 1698431365
transform 1 0 39312 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_364
timestamp 1698431365
transform 1 0 42112 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_384
timestamp 1698431365
transform 1 0 44352 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_387
timestamp 1698431365
transform 1 0 44688 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_391
timestamp 1698431365
transform 1 0 45136 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_393
timestamp 1698431365
transform 1 0 45360 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_439
timestamp 1698431365
transform 1 0 50512 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_457
timestamp 1698431365
transform 1 0 52528 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_489
timestamp 1698431365
transform 1 0 56112 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_505
timestamp 1698431365
transform 1 0 57904 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_6
timestamp 1698431365
transform 1 0 2016 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_22
timestamp 1698431365
transform 1 0 3808 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_30
timestamp 1698431365
transform 1 0 4704 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_34
timestamp 1698431365
transform 1 0 5152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_36
timestamp 1698431365
transform 1 0 5376 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_47
timestamp 1698431365
transform 1 0 6608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_49
timestamp 1698431365
transform 1 0 6832 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_66
timestamp 1698431365
transform 1 0 8736 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_76
timestamp 1698431365
transform 1 0 9856 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_96
timestamp 1698431365
transform 1 0 12096 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_98
timestamp 1698431365
transform 1 0 12320 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_101
timestamp 1698431365
transform 1 0 12656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698431365
transform 1 0 16912 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_144
timestamp 1698431365
transform 1 0 17472 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_161
timestamp 1698431365
transform 1 0 19376 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_163
timestamp 1698431365
transform 1 0 19600 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_189
timestamp 1698431365
transform 1 0 22512 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_225
timestamp 1698431365
transform 1 0 26544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_229
timestamp 1698431365
transform 1 0 26992 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_233
timestamp 1698431365
transform 1 0 27440 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_235
timestamp 1698431365
transform 1 0 27664 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_238
timestamp 1698431365
transform 1 0 28000 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_268
timestamp 1698431365
transform 1 0 31360 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_272
timestamp 1698431365
transform 1 0 31808 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_344
timestamp 1698431365
transform 1 0 39872 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_348
timestamp 1698431365
transform 1 0 40320 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_352
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_356
timestamp 1698431365
transform 1 0 41216 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_377
timestamp 1698431365
transform 1 0 43568 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_409
timestamp 1698431365
transform 1 0 47152 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_417
timestamp 1698431365
transform 1 0 48048 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_419
timestamp 1698431365
transform 1 0 48272 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_422
timestamp 1698431365
transform 1 0 48608 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_426
timestamp 1698431365
transform 1 0 49056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_446
timestamp 1698431365
transform 1 0 51296 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_478
timestamp 1698431365
transform 1 0 54880 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_486
timestamp 1698431365
transform 1 0 55776 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_492
timestamp 1698431365
transform 1 0 56448 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_500
timestamp 1698431365
transform 1 0 57344 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_504
timestamp 1698431365
transform 1 0 57792 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_57
timestamp 1698431365
transform 1 0 7728 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_73
timestamp 1698431365
transform 1 0 9520 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_77
timestamp 1698431365
transform 1 0 9968 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_102
timestamp 1698431365
transform 1 0 12768 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_104
timestamp 1698431365
transform 1 0 12992 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_139
timestamp 1698431365
transform 1 0 16912 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_171
timestamp 1698431365
transform 1 0 20496 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_213
timestamp 1698431365
transform 1 0 25200 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_236
timestamp 1698431365
transform 1 0 27776 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_251
timestamp 1698431365
transform 1 0 29456 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_267
timestamp 1698431365
transform 1 0 31248 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_327
timestamp 1698431365
transform 1 0 37968 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_329
timestamp 1698431365
transform 1 0 38192 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_352
timestamp 1698431365
transform 1 0 40768 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_384
timestamp 1698431365
transform 1 0 44352 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_387
timestamp 1698431365
transform 1 0 44688 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_404
timestamp 1698431365
transform 1 0 46592 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_420
timestamp 1698431365
transform 1 0 48384 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_432
timestamp 1698431365
transform 1 0 49728 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_448
timestamp 1698431365
transform 1 0 51520 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_452
timestamp 1698431365
transform 1 0 51968 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_454
timestamp 1698431365
transform 1 0 52192 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_457
timestamp 1698431365
transform 1 0 52528 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_473
timestamp 1698431365
transform 1 0 54320 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_481
timestamp 1698431365
transform 1 0 55216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_18
timestamp 1698431365
transform 1 0 3360 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_26
timestamp 1698431365
transform 1 0 4256 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_30
timestamp 1698431365
transform 1 0 4704 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_49
timestamp 1698431365
transform 1 0 6832 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_51
timestamp 1698431365
transform 1 0 7056 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_76
timestamp 1698431365
transform 1 0 9856 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_94
timestamp 1698431365
transform 1 0 11872 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_96
timestamp 1698431365
transform 1 0 12096 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_126
timestamp 1698431365
transform 1 0 15456 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_130
timestamp 1698431365
transform 1 0 15904 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_134
timestamp 1698431365
transform 1 0 16352 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_138
timestamp 1698431365
transform 1 0 16800 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_144
timestamp 1698431365
transform 1 0 17472 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_270
timestamp 1698431365
transform 1 0 31584 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_292
timestamp 1698431365
transform 1 0 34048 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_309
timestamp 1698431365
transform 1 0 35952 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_325
timestamp 1698431365
transform 1 0 37744 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_329
timestamp 1698431365
transform 1 0 38192 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_345
timestamp 1698431365
transform 1 0 39984 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_349
timestamp 1698431365
transform 1 0 40432 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_358
timestamp 1698431365
transform 1 0 41440 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_375
timestamp 1698431365
transform 1 0 43344 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_383
timestamp 1698431365
transform 1 0 44240 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_385
timestamp 1698431365
transform 1 0 44464 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_408
timestamp 1698431365
transform 1 0 47040 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_416
timestamp 1698431365
transform 1 0 47936 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_434
timestamp 1698431365
transform 1 0 49952 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_466
timestamp 1698431365
transform 1 0 53536 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_482
timestamp 1698431365
transform 1 0 55328 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_492
timestamp 1698431365
transform 1 0 56448 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_508
timestamp 1698431365
transform 1 0 58240 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_41
timestamp 1698431365
transform 1 0 5936 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_111
timestamp 1698431365
transform 1 0 13776 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_133
timestamp 1698431365
transform 1 0 16240 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_135
timestamp 1698431365
transform 1 0 16464 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_168
timestamp 1698431365
transform 1 0 20160 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_172
timestamp 1698431365
transform 1 0 20608 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_227
timestamp 1698431365
transform 1 0 26768 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_235
timestamp 1698431365
transform 1 0 27664 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_255
timestamp 1698431365
transform 1 0 29904 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_263
timestamp 1698431365
transform 1 0 30800 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_304
timestamp 1698431365
transform 1 0 35392 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_312
timestamp 1698431365
transform 1 0 36288 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_314
timestamp 1698431365
transform 1 0 36512 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_349
timestamp 1698431365
transform 1 0 40432 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_370
timestamp 1698431365
transform 1 0 42784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_387
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_391
timestamp 1698431365
transform 1 0 45136 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_400
timestamp 1698431365
transform 1 0 46144 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_417
timestamp 1698431365
transform 1 0 48048 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_425
timestamp 1698431365
transform 1 0 48944 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_429
timestamp 1698431365
transform 1 0 49392 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_437
timestamp 1698431365
transform 1 0 50288 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_453
timestamp 1698431365
transform 1 0 52080 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_457
timestamp 1698431365
transform 1 0 52528 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_473
timestamp 1698431365
transform 1 0 54320 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_481
timestamp 1698431365
transform 1 0 55216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_6
timestamp 1698431365
transform 1 0 2016 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_38
timestamp 1698431365
transform 1 0 5600 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_40
timestamp 1698431365
transform 1 0 5824 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_49
timestamp 1698431365
transform 1 0 6832 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_61
timestamp 1698431365
transform 1 0 8176 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_90
timestamp 1698431365
transform 1 0 11424 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698431365
transform 1 0 16912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_200
timestamp 1698431365
transform 1 0 23744 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_251
timestamp 1698431365
transform 1 0 29456 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_255
timestamp 1698431365
transform 1 0 29904 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_259
timestamp 1698431365
transform 1 0 30352 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_273
timestamp 1698431365
transform 1 0 31920 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_277
timestamp 1698431365
transform 1 0 32368 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698431365
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_288
timestamp 1698431365
transform 1 0 33600 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_296
timestamp 1698431365
transform 1 0 34496 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_298
timestamp 1698431365
transform 1 0 34720 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_312
timestamp 1698431365
transform 1 0 36288 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_314
timestamp 1698431365
transform 1 0 36512 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_323
timestamp 1698431365
transform 1 0 37520 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_338
timestamp 1698431365
transform 1 0 39200 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_346
timestamp 1698431365
transform 1 0 40096 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_352
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_378
timestamp 1698431365
transform 1 0 43680 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_394
timestamp 1698431365
transform 1 0 45472 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_408
timestamp 1698431365
transform 1 0 47040 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_416
timestamp 1698431365
transform 1 0 47936 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_422
timestamp 1698431365
transform 1 0 48608 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_486
timestamp 1698431365
transform 1 0 55776 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_492
timestamp 1698431365
transform 1 0 56448 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_508
timestamp 1698431365
transform 1 0 58240 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_43
timestamp 1698431365
transform 1 0 6160 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_47
timestamp 1698431365
transform 1 0 6608 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_56
timestamp 1698431365
transform 1 0 7616 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_64
timestamp 1698431365
transform 1 0 8512 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_66
timestamp 1698431365
transform 1 0 8736 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_92
timestamp 1698431365
transform 1 0 11648 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_153
timestamp 1698431365
transform 1 0 18480 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_155
timestamp 1698431365
transform 1 0 18704 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_172
timestamp 1698431365
transform 1 0 20608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698431365
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_197
timestamp 1698431365
transform 1 0 23408 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_199
timestamp 1698431365
transform 1 0 23632 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_260
timestamp 1698431365
transform 1 0 30464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_264
timestamp 1698431365
transform 1 0 30912 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_266
timestamp 1698431365
transform 1 0 31136 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_277
timestamp 1698431365
transform 1 0 32368 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_285
timestamp 1698431365
transform 1 0 33264 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_289
timestamp 1698431365
transform 1 0 33712 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_313
timestamp 1698431365
transform 1 0 36400 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_335
timestamp 1698431365
transform 1 0 38864 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_351
timestamp 1698431365
transform 1 0 40656 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_359
timestamp 1698431365
transform 1 0 41552 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_363
timestamp 1698431365
transform 1 0 42000 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_365
timestamp 1698431365
transform 1 0 42224 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_378
timestamp 1698431365
transform 1 0 43680 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_382
timestamp 1698431365
transform 1 0 44128 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_384
timestamp 1698431365
transform 1 0 44352 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_387
timestamp 1698431365
transform 1 0 44688 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_403
timestamp 1698431365
transform 1 0 46480 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_410
timestamp 1698431365
transform 1 0 47264 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_442
timestamp 1698431365
transform 1 0 50848 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_450
timestamp 1698431365
transform 1 0 51744 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_454
timestamp 1698431365
transform 1 0 52192 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_457
timestamp 1698431365
transform 1 0 52528 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_473
timestamp 1698431365
transform 1 0 54320 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_481
timestamp 1698431365
transform 1 0 55216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_10
timestamp 1698431365
transform 1 0 2464 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_26
timestamp 1698431365
transform 1 0 4256 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_28
timestamp 1698431365
transform 1 0 4480 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_52
timestamp 1698431365
transform 1 0 7168 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_56
timestamp 1698431365
transform 1 0 7616 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_58
timestamp 1698431365
transform 1 0 7840 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_67
timestamp 1698431365
transform 1 0 8848 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_69
timestamp 1698431365
transform 1 0 9072 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_74
timestamp 1698431365
transform 1 0 9632 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_103
timestamp 1698431365
transform 1 0 12880 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_136
timestamp 1698431365
transform 1 0 16576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_144
timestamp 1698431365
transform 1 0 17472 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_197
timestamp 1698431365
transform 1 0 23408 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_208
timestamp 1698431365
transform 1 0 24640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_245
timestamp 1698431365
transform 1 0 28784 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_314
timestamp 1698431365
transform 1 0 36512 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_330
timestamp 1698431365
transform 1 0 38304 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_340
timestamp 1698431365
transform 1 0 39424 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_344
timestamp 1698431365
transform 1 0 39872 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_348
timestamp 1698431365
transform 1 0 40320 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_352
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_360
timestamp 1698431365
transform 1 0 41664 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_364
timestamp 1698431365
transform 1 0 42112 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_399
timestamp 1698431365
transform 1 0 46032 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_415
timestamp 1698431365
transform 1 0 47824 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_419
timestamp 1698431365
transform 1 0 48272 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_422
timestamp 1698431365
transform 1 0 48608 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_486
timestamp 1698431365
transform 1 0 55776 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_492
timestamp 1698431365
transform 1 0 56448 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_500
timestamp 1698431365
transform 1 0 57344 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_504
timestamp 1698431365
transform 1 0 57792 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_28
timestamp 1698431365
transform 1 0 4480 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_32
timestamp 1698431365
transform 1 0 4928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_75
timestamp 1698431365
transform 1 0 9744 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_79
timestamp 1698431365
transform 1 0 10192 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_98
timestamp 1698431365
transform 1 0 12320 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_102
timestamp 1698431365
transform 1 0 12768 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_115
timestamp 1698431365
transform 1 0 14224 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_124
timestamp 1698431365
transform 1 0 15232 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_138
timestamp 1698431365
transform 1 0 16800 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_158
timestamp 1698431365
transform 1 0 19040 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_160
timestamp 1698431365
transform 1 0 19264 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_163
timestamp 1698431365
transform 1 0 19600 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_167
timestamp 1698431365
transform 1 0 20048 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_171
timestamp 1698431365
transform 1 0 20496 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_185
timestamp 1698431365
transform 1 0 22064 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_189
timestamp 1698431365
transform 1 0 22512 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_264
timestamp 1698431365
transform 1 0 30912 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_305
timestamp 1698431365
transform 1 0 35504 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_309
timestamp 1698431365
transform 1 0 35952 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_313
timestamp 1698431365
transform 1 0 36400 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_325
timestamp 1698431365
transform 1 0 37744 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_329
timestamp 1698431365
transform 1 0 38192 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_331
timestamp 1698431365
transform 1 0 38416 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_374
timestamp 1698431365
transform 1 0 43232 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_378
timestamp 1698431365
transform 1 0 43680 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_382
timestamp 1698431365
transform 1 0 44128 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_384
timestamp 1698431365
transform 1 0 44352 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_387
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_451
timestamp 1698431365
transform 1 0 51856 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_457
timestamp 1698431365
transform 1 0 52528 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_489
timestamp 1698431365
transform 1 0 56112 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_18
timestamp 1698431365
transform 1 0 3360 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_26
timestamp 1698431365
transform 1 0 4256 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_65
timestamp 1698431365
transform 1 0 8624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_69
timestamp 1698431365
transform 1 0 9072 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_78
timestamp 1698431365
transform 1 0 10080 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_80
timestamp 1698431365
transform 1 0 10304 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_103
timestamp 1698431365
transform 1 0 12880 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_119
timestamp 1698431365
transform 1 0 14672 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_129
timestamp 1698431365
transform 1 0 15792 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_131
timestamp 1698431365
transform 1 0 16016 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_150
timestamp 1698431365
transform 1 0 18144 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_159
timestamp 1698431365
transform 1 0 19152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_163
timestamp 1698431365
transform 1 0 19600 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_167
timestamp 1698431365
transform 1 0 20048 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_183
timestamp 1698431365
transform 1 0 21840 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_191
timestamp 1698431365
transform 1 0 22736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_195
timestamp 1698431365
transform 1 0 23184 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_204
timestamp 1698431365
transform 1 0 24192 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_226
timestamp 1698431365
transform 1 0 26656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_230
timestamp 1698431365
transform 1 0 27104 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_234
timestamp 1698431365
transform 1 0 27552 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_245
timestamp 1698431365
transform 1 0 28784 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_249
timestamp 1698431365
transform 1 0 29232 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_253
timestamp 1698431365
transform 1 0 29680 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_256
timestamp 1698431365
transform 1 0 30016 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_260
timestamp 1698431365
transform 1 0 30464 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_262
timestamp 1698431365
transform 1 0 30688 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_265
timestamp 1698431365
transform 1 0 31024 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_273
timestamp 1698431365
transform 1 0 31920 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_277
timestamp 1698431365
transform 1 0 32368 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_298
timestamp 1698431365
transform 1 0 34720 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_302
timestamp 1698431365
transform 1 0 35168 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_335
timestamp 1698431365
transform 1 0 38864 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_343
timestamp 1698431365
transform 1 0 39760 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_347
timestamp 1698431365
transform 1 0 40208 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_349
timestamp 1698431365
transform 1 0 40432 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_386
timestamp 1698431365
transform 1 0 44576 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_418
timestamp 1698431365
transform 1 0 48160 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_422
timestamp 1698431365
transform 1 0 48608 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_486
timestamp 1698431365
transform 1 0 55776 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_492
timestamp 1698431365
transform 1 0 56448 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_508
timestamp 1698431365
transform 1 0 58240 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_28
timestamp 1698431365
transform 1 0 4480 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_32
timestamp 1698431365
transform 1 0 4928 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_45
timestamp 1698431365
transform 1 0 6384 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_55
timestamp 1698431365
transform 1 0 7504 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_63
timestamp 1698431365
transform 1 0 8400 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_67
timestamp 1698431365
transform 1 0 8848 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_85
timestamp 1698431365
transform 1 0 10864 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_89
timestamp 1698431365
transform 1 0 11312 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_98
timestamp 1698431365
transform 1 0 12320 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_102
timestamp 1698431365
transform 1 0 12768 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_139
timestamp 1698431365
transform 1 0 16912 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_143
timestamp 1698431365
transform 1 0 17360 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_152
timestamp 1698431365
transform 1 0 18368 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_156
timestamp 1698431365
transform 1 0 18816 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_162
timestamp 1698431365
transform 1 0 19488 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_166
timestamp 1698431365
transform 1 0 19936 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_185
timestamp 1698431365
transform 1 0 22064 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_189
timestamp 1698431365
transform 1 0 22512 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_193
timestamp 1698431365
transform 1 0 22960 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_201
timestamp 1698431365
transform 1 0 23856 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_203
timestamp 1698431365
transform 1 0 24080 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_223
timestamp 1698431365
transform 1 0 26320 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_239
timestamp 1698431365
transform 1 0 28112 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_243
timestamp 1698431365
transform 1 0 28560 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_253
timestamp 1698431365
transform 1 0 29680 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_261
timestamp 1698431365
transform 1 0 30576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_278
timestamp 1698431365
transform 1 0 32480 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_280
timestamp 1698431365
transform 1 0 32704 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_289
timestamp 1698431365
transform 1 0 33712 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_293
timestamp 1698431365
transform 1 0 34160 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_309
timestamp 1698431365
transform 1 0 35952 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_313
timestamp 1698431365
transform 1 0 36400 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_326
timestamp 1698431365
transform 1 0 37856 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_334
timestamp 1698431365
transform 1 0 38752 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_366
timestamp 1698431365
transform 1 0 42336 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_382
timestamp 1698431365
transform 1 0 44128 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_384
timestamp 1698431365
transform 1 0 44352 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_387
timestamp 1698431365
transform 1 0 44688 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_451
timestamp 1698431365
transform 1 0 51856 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_457
timestamp 1698431365
transform 1 0 52528 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_489
timestamp 1698431365
transform 1 0 56112 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_28
timestamp 1698431365
transform 1 0 4480 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_60
timestamp 1698431365
transform 1 0 8064 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_68
timestamp 1698431365
transform 1 0 8960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_74
timestamp 1698431365
transform 1 0 9632 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_89
timestamp 1698431365
transform 1 0 11312 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_105
timestamp 1698431365
transform 1 0 13104 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_111
timestamp 1698431365
transform 1 0 13776 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_118
timestamp 1698431365
transform 1 0 14560 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_122
timestamp 1698431365
transform 1 0 15008 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_134
timestamp 1698431365
transform 1 0 16352 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_138
timestamp 1698431365
transform 1 0 16800 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_161
timestamp 1698431365
transform 1 0 19376 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_169
timestamp 1698431365
transform 1 0 20272 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_190
timestamp 1698431365
transform 1 0 22624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_194
timestamp 1698431365
transform 1 0 23072 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_202
timestamp 1698431365
transform 1 0 23968 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_206
timestamp 1698431365
transform 1 0 24416 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_220
timestamp 1698431365
transform 1 0 25984 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_224
timestamp 1698431365
transform 1 0 26432 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_232
timestamp 1698431365
transform 1 0 27328 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_236
timestamp 1698431365
transform 1 0 27776 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698431365
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_318
timestamp 1698431365
transform 1 0 36960 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_328
timestamp 1698431365
transform 1 0 38080 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_345
timestamp 1698431365
transform 1 0 39984 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_349
timestamp 1698431365
transform 1 0 40432 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_352
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_368
timestamp 1698431365
transform 1 0 42560 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_403
timestamp 1698431365
transform 1 0 46480 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_419
timestamp 1698431365
transform 1 0 48272 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_422
timestamp 1698431365
transform 1 0 48608 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_486
timestamp 1698431365
transform 1 0 55776 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_492
timestamp 1698431365
transform 1 0 56448 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_508
timestamp 1698431365
transform 1 0 58240 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_28
timestamp 1698431365
transform 1 0 4480 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_32
timestamp 1698431365
transform 1 0 4928 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_43
timestamp 1698431365
transform 1 0 6160 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_51
timestamp 1698431365
transform 1 0 7056 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_55
timestamp 1698431365
transform 1 0 7504 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_91
timestamp 1698431365
transform 1 0 11536 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_95
timestamp 1698431365
transform 1 0 11984 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_103
timestamp 1698431365
transform 1 0 12880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_114
timestamp 1698431365
transform 1 0 14112 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_130
timestamp 1698431365
transform 1 0 15904 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_155
timestamp 1698431365
transform 1 0 18704 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_157
timestamp 1698431365
transform 1 0 18928 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_172
timestamp 1698431365
transform 1 0 20608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_174
timestamp 1698431365
transform 1 0 20832 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_186
timestamp 1698431365
transform 1 0 22176 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_190
timestamp 1698431365
transform 1 0 22624 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_198
timestamp 1698431365
transform 1 0 23520 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_255
timestamp 1698431365
transform 1 0 29904 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_259
timestamp 1698431365
transform 1 0 30352 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_267
timestamp 1698431365
transform 1 0 31248 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_289
timestamp 1698431365
transform 1 0 33712 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_293
timestamp 1698431365
transform 1 0 34160 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_309
timestamp 1698431365
transform 1 0 35952 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_313
timestamp 1698431365
transform 1 0 36400 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_319
timestamp 1698431365
transform 1 0 37072 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_326
timestamp 1698431365
transform 1 0 37856 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_330
timestamp 1698431365
transform 1 0 38304 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_365
timestamp 1698431365
transform 1 0 42224 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_373
timestamp 1698431365
transform 1 0 43120 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_377
timestamp 1698431365
transform 1 0 43568 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_379
timestamp 1698431365
transform 1 0 43792 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_387
timestamp 1698431365
transform 1 0 44688 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_400
timestamp 1698431365
transform 1 0 46144 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_432
timestamp 1698431365
transform 1 0 49728 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_448
timestamp 1698431365
transform 1 0 51520 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_452
timestamp 1698431365
transform 1 0 51968 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_454
timestamp 1698431365
transform 1 0 52192 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_457
timestamp 1698431365
transform 1 0 52528 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_489
timestamp 1698431365
transform 1 0 56112 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_505
timestamp 1698431365
transform 1 0 57904 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_28
timestamp 1698431365
transform 1 0 4480 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_64
timestamp 1698431365
transform 1 0 8512 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_68
timestamp 1698431365
transform 1 0 8960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_78
timestamp 1698431365
transform 1 0 10080 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_94
timestamp 1698431365
transform 1 0 11872 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_98
timestamp 1698431365
transform 1 0 12320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_133
timestamp 1698431365
transform 1 0 16240 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_137
timestamp 1698431365
transform 1 0 16688 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_139
timestamp 1698431365
transform 1 0 16912 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_149
timestamp 1698431365
transform 1 0 18032 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_155
timestamp 1698431365
transform 1 0 18704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_209
timestamp 1698431365
transform 1 0 24752 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_220
timestamp 1698431365
transform 1 0 25984 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_224
timestamp 1698431365
transform 1 0 26432 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698431365
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_292
timestamp 1698431365
transform 1 0 34048 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_324
timestamp 1698431365
transform 1 0 37632 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_328
timestamp 1698431365
transform 1 0 38080 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_330
timestamp 1698431365
transform 1 0 38304 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_345
timestamp 1698431365
transform 1 0 39984 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_349
timestamp 1698431365
transform 1 0 40432 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_365
timestamp 1698431365
transform 1 0 42224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_401
timestamp 1698431365
transform 1 0 46256 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_412
timestamp 1698431365
transform 1 0 47488 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_422
timestamp 1698431365
transform 1 0 48608 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_486
timestamp 1698431365
transform 1 0 55776 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_492
timestamp 1698431365
transform 1 0 56448 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_500
timestamp 1698431365
transform 1 0 57344 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_12
timestamp 1698431365
transform 1 0 2688 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_30
timestamp 1698431365
transform 1 0 4704 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698431365
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_139
timestamp 1698431365
transform 1 0 16912 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_147
timestamp 1698431365
transform 1 0 17808 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_155
timestamp 1698431365
transform 1 0 18704 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_162
timestamp 1698431365
transform 1 0 19488 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_170
timestamp 1698431365
transform 1 0 20384 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_174
timestamp 1698431365
transform 1 0 20832 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_213
timestamp 1698431365
transform 1 0 25200 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_217
timestamp 1698431365
transform 1 0 25648 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_221
timestamp 1698431365
transform 1 0 26096 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_237
timestamp 1698431365
transform 1 0 27888 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_251
timestamp 1698431365
transform 1 0 29456 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_253
timestamp 1698431365
transform 1 0 29680 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_288
timestamp 1698431365
transform 1 0 33600 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_297
timestamp 1698431365
transform 1 0 34608 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_313
timestamp 1698431365
transform 1 0 36400 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_321
timestamp 1698431365
transform 1 0 37296 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_341
timestamp 1698431365
transform 1 0 39536 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_373
timestamp 1698431365
transform 1 0 43120 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_381
timestamp 1698431365
transform 1 0 44016 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_387
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_395
timestamp 1698431365
transform 1 0 45584 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_399
timestamp 1698431365
transform 1 0 46032 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_402
timestamp 1698431365
transform 1 0 46368 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_418
timestamp 1698431365
transform 1 0 48160 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_420
timestamp 1698431365
transform 1 0 48384 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_429
timestamp 1698431365
transform 1 0 49392 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_445
timestamp 1698431365
transform 1 0 51184 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_453
timestamp 1698431365
transform 1 0 52080 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_457
timestamp 1698431365
transform 1 0 52528 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_489
timestamp 1698431365
transform 1 0 56112 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_505
timestamp 1698431365
transform 1 0 57904 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_6
timestamp 1698431365
transform 1 0 2016 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_88
timestamp 1698431365
transform 1 0 11200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_158
timestamp 1698431365
transform 1 0 19040 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_162
timestamp 1698431365
transform 1 0 19488 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_168
timestamp 1698431365
transform 1 0 20160 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_172
timestamp 1698431365
transform 1 0 20608 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_188
timestamp 1698431365
transform 1 0 22400 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_200
timestamp 1698431365
transform 1 0 23744 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_219
timestamp 1698431365
transform 1 0 25872 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_263
timestamp 1698431365
transform 1 0 30800 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_279
timestamp 1698431365
transform 1 0 32592 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_286
timestamp 1698431365
transform 1 0 33376 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_333
timestamp 1698431365
transform 1 0 38640 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_349
timestamp 1698431365
transform 1 0 40432 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_368
timestamp 1698431365
transform 1 0 42560 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_372
timestamp 1698431365
transform 1 0 43008 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_375
timestamp 1698431365
transform 1 0 43344 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_381
timestamp 1698431365
transform 1 0 44016 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_397
timestamp 1698431365
transform 1 0 45808 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_405
timestamp 1698431365
transform 1 0 46704 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_414
timestamp 1698431365
transform 1 0 47712 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_422
timestamp 1698431365
transform 1 0 48608 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_426
timestamp 1698431365
transform 1 0 49056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_428
timestamp 1698431365
transform 1 0 49280 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_439
timestamp 1698431365
transform 1 0 50512 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_471
timestamp 1698431365
transform 1 0 54096 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_487
timestamp 1698431365
transform 1 0 55888 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_489
timestamp 1698431365
transform 1 0 56112 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_492
timestamp 1698431365
transform 1 0 56448 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_508
timestamp 1698431365
transform 1 0 58240 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_8
timestamp 1698431365
transform 1 0 2240 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_12
timestamp 1698431365
transform 1 0 2688 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_28
timestamp 1698431365
transform 1 0 4480 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_32
timestamp 1698431365
transform 1 0 4928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_53
timestamp 1698431365
transform 1 0 7280 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_61
timestamp 1698431365
transform 1 0 8176 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_98
timestamp 1698431365
transform 1 0 12320 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_102
timestamp 1698431365
transform 1 0 12768 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_104
timestamp 1698431365
transform 1 0 12992 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_147
timestamp 1698431365
transform 1 0 17808 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_151
timestamp 1698431365
transform 1 0 18256 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_172
timestamp 1698431365
transform 1 0 20608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_174
timestamp 1698431365
transform 1 0 20832 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_181
timestamp 1698431365
transform 1 0 21616 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_191
timestamp 1698431365
transform 1 0 22736 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_195
timestamp 1698431365
transform 1 0 23184 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_197
timestamp 1698431365
transform 1 0 23408 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_200
timestamp 1698431365
transform 1 0 23744 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_231
timestamp 1698431365
transform 1 0 27216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_235
timestamp 1698431365
transform 1 0 27664 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_249
timestamp 1698431365
transform 1 0 29232 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_256
timestamp 1698431365
transform 1 0 30016 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_260
timestamp 1698431365
transform 1 0 30464 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_292
timestamp 1698431365
transform 1 0 34048 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_295
timestamp 1698431365
transform 1 0 34384 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_303
timestamp 1698431365
transform 1 0 35280 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_307
timestamp 1698431365
transform 1 0 35728 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_321
timestamp 1698431365
transform 1 0 37296 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_356
timestamp 1698431365
transform 1 0 41216 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_360
timestamp 1698431365
transform 1 0 41664 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_362
timestamp 1698431365
transform 1 0 41888 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_381
timestamp 1698431365
transform 1 0 44016 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_416
timestamp 1698431365
transform 1 0 47936 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_437
timestamp 1698431365
transform 1 0 50288 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_450
timestamp 1698431365
transform 1 0 51744 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_454
timestamp 1698431365
transform 1 0 52192 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_475
timestamp 1698431365
transform 1 0 54544 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_34
timestamp 1698431365
transform 1 0 5152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_80
timestamp 1698431365
transform 1 0 10304 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_122
timestamp 1698431365
transform 1 0 15008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_126
timestamp 1698431365
transform 1 0 15456 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_134
timestamp 1698431365
transform 1 0 16352 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_150
timestamp 1698431365
transform 1 0 18144 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_170
timestamp 1698431365
transform 1 0 20384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_172
timestamp 1698431365
transform 1 0 20608 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_185
timestamp 1698431365
transform 1 0 22064 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_189
timestamp 1698431365
transform 1 0 22512 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_193
timestamp 1698431365
transform 1 0 22960 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_200
timestamp 1698431365
transform 1 0 23744 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_208
timestamp 1698431365
transform 1 0 24640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_214
timestamp 1698431365
transform 1 0 25312 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_225
timestamp 1698431365
transform 1 0 26544 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_241
timestamp 1698431365
transform 1 0 28336 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_245
timestamp 1698431365
transform 1 0 28784 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_268
timestamp 1698431365
transform 1 0 31360 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698431365
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_286
timestamp 1698431365
transform 1 0 33376 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_343
timestamp 1698431365
transform 1 0 39760 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_386
timestamp 1698431365
transform 1 0 44576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_388
timestamp 1698431365
transform 1 0 44800 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_395
timestamp 1698431365
transform 1 0 45584 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_410
timestamp 1698431365
transform 1 0 47264 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_418
timestamp 1698431365
transform 1 0 48160 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_422
timestamp 1698431365
transform 1 0 48608 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_430
timestamp 1698431365
transform 1 0 49504 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_445
timestamp 1698431365
transform 1 0 51184 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_449
timestamp 1698431365
transform 1 0 51632 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_477
timestamp 1698431365
transform 1 0 54768 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_479
timestamp 1698431365
transform 1 0 54992 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_486
timestamp 1698431365
transform 1 0 55776 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_492
timestamp 1698431365
transform 1 0 56448 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_508
timestamp 1698431365
transform 1 0 58240 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_83
timestamp 1698431365
transform 1 0 10640 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_87
timestamp 1698431365
transform 1 0 11088 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_91
timestamp 1698431365
transform 1 0 11536 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_99
timestamp 1698431365
transform 1 0 12432 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_113
timestamp 1698431365
transform 1 0 14000 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_117
timestamp 1698431365
transform 1 0 14448 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_124
timestamp 1698431365
transform 1 0 15232 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_140
timestamp 1698431365
transform 1 0 17024 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_148
timestamp 1698431365
transform 1 0 17920 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_157
timestamp 1698431365
transform 1 0 18928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_159
timestamp 1698431365
transform 1 0 19152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_170
timestamp 1698431365
transform 1 0 20384 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_174
timestamp 1698431365
transform 1 0 20832 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_195
timestamp 1698431365
transform 1 0 23184 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_211
timestamp 1698431365
transform 1 0 24976 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_221
timestamp 1698431365
transform 1 0 26096 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_234
timestamp 1698431365
transform 1 0 27552 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_242
timestamp 1698431365
transform 1 0 28448 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_253
timestamp 1698431365
transform 1 0 29680 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_283
timestamp 1698431365
transform 1 0 33040 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_295
timestamp 1698431365
transform 1 0 34384 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698431365
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_342
timestamp 1698431365
transform 1 0 39648 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_352
timestamp 1698431365
transform 1 0 40768 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_368
timestamp 1698431365
transform 1 0 42560 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_372
timestamp 1698431365
transform 1 0 43008 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_379
timestamp 1698431365
transform 1 0 43792 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_383
timestamp 1698431365
transform 1 0 44240 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_392
timestamp 1698431365
transform 1 0 45248 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_400
timestamp 1698431365
transform 1 0 46144 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_407
timestamp 1698431365
transform 1 0 46928 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_435
timestamp 1698431365
transform 1 0 50064 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_439
timestamp 1698431365
transform 1 0 50512 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_494
timestamp 1698431365
transform 1 0 56672 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_502
timestamp 1698431365
transform 1 0 57568 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_506
timestamp 1698431365
transform 1 0 58016 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_508
timestamp 1698431365
transform 1 0 58240 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_28
timestamp 1698431365
transform 1 0 4480 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_44
timestamp 1698431365
transform 1 0 6272 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_56
timestamp 1698431365
transform 1 0 7616 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698431365
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_85
timestamp 1698431365
transform 1 0 10864 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_102
timestamp 1698431365
transform 1 0 12768 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_104
timestamp 1698431365
transform 1 0 12992 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_135
timestamp 1698431365
transform 1 0 16464 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_139
timestamp 1698431365
transform 1 0 16912 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_150
timestamp 1698431365
transform 1 0 18144 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_160
timestamp 1698431365
transform 1 0 19264 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_172
timestamp 1698431365
transform 1 0 20608 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_176
timestamp 1698431365
transform 1 0 21056 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_180
timestamp 1698431365
transform 1 0 21504 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_188
timestamp 1698431365
transform 1 0 22400 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_192
timestamp 1698431365
transform 1 0 22848 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_217
timestamp 1698431365
transform 1 0 25648 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_219
timestamp 1698431365
transform 1 0 25872 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_222
timestamp 1698431365
transform 1 0 26208 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_226
timestamp 1698431365
transform 1 0 26656 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_232
timestamp 1698431365
transform 1 0 27328 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_240
timestamp 1698431365
transform 1 0 28224 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_243
timestamp 1698431365
transform 1 0 28560 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_247
timestamp 1698431365
transform 1 0 29008 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_262
timestamp 1698431365
transform 1 0 30688 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_297
timestamp 1698431365
transform 1 0 34608 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_309
timestamp 1698431365
transform 1 0 35952 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_314
timestamp 1698431365
transform 1 0 36512 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_318
timestamp 1698431365
transform 1 0 36960 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_325
timestamp 1698431365
transform 1 0 37744 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_342
timestamp 1698431365
transform 1 0 39648 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_354
timestamp 1698431365
transform 1 0 40992 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_360
timestamp 1698431365
transform 1 0 41664 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_364
timestamp 1698431365
transform 1 0 42112 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_403
timestamp 1698431365
transform 1 0 46480 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_419
timestamp 1698431365
transform 1 0 48272 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_434
timestamp 1698431365
transform 1 0 49952 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_450
timestamp 1698431365
transform 1 0 51744 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_454
timestamp 1698431365
transform 1 0 52192 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_467
timestamp 1698431365
transform 1 0 53648 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_482
timestamp 1698431365
transform 1 0 55328 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_492
timestamp 1698431365
transform 1 0 56448 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_508
timestamp 1698431365
transform 1 0 58240 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_28
timestamp 1698431365
transform 1 0 4480 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_32
timestamp 1698431365
transform 1 0 4928 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_53
timestamp 1698431365
transform 1 0 7280 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_60
timestamp 1698431365
transform 1 0 8064 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_88
timestamp 1698431365
transform 1 0 11200 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_92
timestamp 1698431365
transform 1 0 11648 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_143
timestamp 1698431365
transform 1 0 17360 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_145
timestamp 1698431365
transform 1 0 17584 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_154
timestamp 1698431365
transform 1 0 18592 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_158
timestamp 1698431365
transform 1 0 19040 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_179
timestamp 1698431365
transform 1 0 21392 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_220
timestamp 1698431365
transform 1 0 25984 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_242
timestamp 1698431365
transform 1 0 28448 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_244
timestamp 1698431365
transform 1 0 28672 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_253
timestamp 1698431365
transform 1 0 29680 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_257
timestamp 1698431365
transform 1 0 30128 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_298
timestamp 1698431365
transform 1 0 34720 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_313
timestamp 1698431365
transform 1 0 36400 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_325
timestamp 1698431365
transform 1 0 37744 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_331
timestamp 1698431365
transform 1 0 38416 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_335
timestamp 1698431365
transform 1 0 38864 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_345
timestamp 1698431365
transform 1 0 39984 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_353
timestamp 1698431365
transform 1 0 40880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_370
timestamp 1698431365
transform 1 0 42784 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_378
timestamp 1698431365
transform 1 0 43680 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_382
timestamp 1698431365
transform 1 0 44128 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_384
timestamp 1698431365
transform 1 0 44352 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_433
timestamp 1698431365
transform 1 0 49840 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_451
timestamp 1698431365
transform 1 0 51856 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_457
timestamp 1698431365
transform 1 0 52528 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_465
timestamp 1698431365
transform 1 0 53424 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_475
timestamp 1698431365
transform 1 0 54544 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_10
timestamp 1698431365
transform 1 0 2464 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_42
timestamp 1698431365
transform 1 0 6048 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_46
timestamp 1698431365
transform 1 0 6496 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_48
timestamp 1698431365
transform 1 0 6720 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_63
timestamp 1698431365
transform 1 0 8400 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_80
timestamp 1698431365
transform 1 0 10304 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_90
timestamp 1698431365
transform 1 0 11424 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_98
timestamp 1698431365
transform 1 0 12320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_115
timestamp 1698431365
transform 1 0 14224 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_119
timestamp 1698431365
transform 1 0 14672 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_121
timestamp 1698431365
transform 1 0 14896 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_133
timestamp 1698431365
transform 1 0 16240 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_137
timestamp 1698431365
transform 1 0 16688 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_139
timestamp 1698431365
transform 1 0 16912 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_142
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_160
timestamp 1698431365
transform 1 0 19264 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_180
timestamp 1698431365
transform 1 0 21504 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_187
timestamp 1698431365
transform 1 0 22288 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_195
timestamp 1698431365
transform 1 0 23184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_199
timestamp 1698431365
transform 1 0 23632 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_208
timestamp 1698431365
transform 1 0 24640 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_212
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698431365
transform 1 0 32592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_288
timestamp 1698431365
transform 1 0 33600 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_352
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_368
timestamp 1698431365
transform 1 0 42560 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_376
timestamp 1698431365
transform 1 0 43456 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_380
timestamp 1698431365
transform 1 0 43904 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_404
timestamp 1698431365
transform 1 0 46592 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_422
timestamp 1698431365
transform 1 0 48608 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_430
timestamp 1698431365
transform 1 0 49504 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_469
timestamp 1698431365
transform 1 0 53872 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_479
timestamp 1698431365
transform 1 0 54992 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_483
timestamp 1698431365
transform 1 0 55440 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_492
timestamp 1698431365
transform 1 0 56448 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_508
timestamp 1698431365
transform 1 0 58240 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698431365
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_69
timestamp 1698431365
transform 1 0 9072 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_77
timestamp 1698431365
transform 1 0 9968 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_84
timestamp 1698431365
transform 1 0 10752 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_100
timestamp 1698431365
transform 1 0 12544 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_104
timestamp 1698431365
transform 1 0 12992 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_115
timestamp 1698431365
transform 1 0 14224 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_125
timestamp 1698431365
transform 1 0 15344 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_142
timestamp 1698431365
transform 1 0 17248 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_162
timestamp 1698431365
transform 1 0 19488 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_166
timestamp 1698431365
transform 1 0 19936 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_185
timestamp 1698431365
transform 1 0 22064 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_193
timestamp 1698431365
transform 1 0 22960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_195
timestamp 1698431365
transform 1 0 23184 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_204
timestamp 1698431365
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_206
timestamp 1698431365
transform 1 0 24416 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_217
timestamp 1698431365
transform 1 0 25648 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_219
timestamp 1698431365
transform 1 0 25872 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_255
timestamp 1698431365
transform 1 0 29904 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_259
timestamp 1698431365
transform 1 0 30352 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_263
timestamp 1698431365
transform 1 0 30800 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_265
timestamp 1698431365
transform 1 0 31024 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_291
timestamp 1698431365
transform 1 0 33936 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_317
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_321
timestamp 1698431365
transform 1 0 37296 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_331
timestamp 1698431365
transform 1 0 38416 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_363
timestamp 1698431365
transform 1 0 42000 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_382
timestamp 1698431365
transform 1 0 44128 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_384
timestamp 1698431365
transform 1 0 44352 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_387
timestamp 1698431365
transform 1 0 44688 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_402
timestamp 1698431365
transform 1 0 46368 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_434
timestamp 1698431365
transform 1 0 49952 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_438
timestamp 1698431365
transform 1 0 50400 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_440
timestamp 1698431365
transform 1 0 50624 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_453
timestamp 1698431365
transform 1 0 52080 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_457
timestamp 1698431365
transform 1 0 52528 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_2
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_34
timestamp 1698431365
transform 1 0 5152 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_50
timestamp 1698431365
transform 1 0 6944 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_54
timestamp 1698431365
transform 1 0 7392 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_61
timestamp 1698431365
transform 1 0 8176 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_65
timestamp 1698431365
transform 1 0 8624 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_69
timestamp 1698431365
transform 1 0 9072 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_80
timestamp 1698431365
transform 1 0 10304 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_82
timestamp 1698431365
transform 1 0 10528 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_115
timestamp 1698431365
transform 1 0 14224 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_126
timestamp 1698431365
transform 1 0 15456 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_130
timestamp 1698431365
transform 1 0 15904 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_155
timestamp 1698431365
transform 1 0 18704 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_169
timestamp 1698431365
transform 1 0 20272 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_177
timestamp 1698431365
transform 1 0 21168 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_181
timestamp 1698431365
transform 1 0 21616 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_195
timestamp 1698431365
transform 1 0 23184 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_199
timestamp 1698431365
transform 1 0 23632 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_228
timestamp 1698431365
transform 1 0 26880 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_232
timestamp 1698431365
transform 1 0 27328 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_266
timestamp 1698431365
transform 1 0 31136 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_268
timestamp 1698431365
transform 1 0 31360 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_282
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_288
timestamp 1698431365
transform 1 0 33600 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_292
timestamp 1698431365
transform 1 0 34048 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_296
timestamp 1698431365
transform 1 0 34496 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_312
timestamp 1698431365
transform 1 0 36288 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_340
timestamp 1698431365
transform 1 0 39424 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_348
timestamp 1698431365
transform 1 0 40320 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_352
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_356
timestamp 1698431365
transform 1 0 41216 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_379
timestamp 1698431365
transform 1 0 43792 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_416
timestamp 1698431365
transform 1 0 47936 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_432
timestamp 1698431365
transform 1 0 49728 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_436
timestamp 1698431365
transform 1 0 50176 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_440
timestamp 1698431365
transform 1 0 50624 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_456
timestamp 1698431365
transform 1 0 52416 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_460
timestamp 1698431365
transform 1 0 52864 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_479
timestamp 1698431365
transform 1 0 54992 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_487
timestamp 1698431365
transform 1 0 55888 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_489
timestamp 1698431365
transform 1 0 56112 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_492
timestamp 1698431365
transform 1 0 56448 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_508
timestamp 1698431365
transform 1 0 58240 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_6
timestamp 1698431365
transform 1 0 2016 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_22
timestamp 1698431365
transform 1 0 3808 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_30
timestamp 1698431365
transform 1 0 4704 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698431365
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_78
timestamp 1698431365
transform 1 0 10080 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_80
timestamp 1698431365
transform 1 0 10304 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_115
timestamp 1698431365
transform 1 0 14224 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_129
timestamp 1698431365
transform 1 0 15792 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_133
timestamp 1698431365
transform 1 0 16240 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_171
timestamp 1698431365
transform 1 0 20496 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_192
timestamp 1698431365
transform 1 0 22848 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_201
timestamp 1698431365
transform 1 0 23856 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_203
timestamp 1698431365
transform 1 0 24080 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_214
timestamp 1698431365
transform 1 0 25312 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_218
timestamp 1698431365
transform 1 0 25760 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_222
timestamp 1698431365
transform 1 0 26208 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_244
timestamp 1698431365
transform 1 0 28672 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_255
timestamp 1698431365
transform 1 0 29904 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_263
timestamp 1698431365
transform 1 0 30800 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_267
timestamp 1698431365
transform 1 0 31248 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_269
timestamp 1698431365
transform 1 0 31472 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_296
timestamp 1698431365
transform 1 0 34496 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_312
timestamp 1698431365
transform 1 0 36288 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_314
timestamp 1698431365
transform 1 0 36512 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_317
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_321
timestamp 1698431365
transform 1 0 37296 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_323
timestamp 1698431365
transform 1 0 37520 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_334
timestamp 1698431365
transform 1 0 38752 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_338
timestamp 1698431365
transform 1 0 39200 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_346
timestamp 1698431365
transform 1 0 40096 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_362
timestamp 1698431365
transform 1 0 41888 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_372
timestamp 1698431365
transform 1 0 43008 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_380
timestamp 1698431365
transform 1 0 43904 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_384
timestamp 1698431365
transform 1 0 44352 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_393
timestamp 1698431365
transform 1 0 45360 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_395
timestamp 1698431365
transform 1 0 45584 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_409
timestamp 1698431365
transform 1 0 47152 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_417
timestamp 1698431365
transform 1 0 48048 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_448
timestamp 1698431365
transform 1 0 51520 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_452
timestamp 1698431365
transform 1 0 51968 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_454
timestamp 1698431365
transform 1 0 52192 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_457
timestamp 1698431365
transform 1 0 52528 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_465
timestamp 1698431365
transform 1 0 53424 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_474
timestamp 1698431365
transform 1 0 54432 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_482
timestamp 1698431365
transform 1 0 55328 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_34
timestamp 1698431365
transform 1 0 5152 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_50
timestamp 1698431365
transform 1 0 6944 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_57
timestamp 1698431365
transform 1 0 7728 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_169
timestamp 1698431365
transform 1 0 20272 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_191
timestamp 1698431365
transform 1 0 22736 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_195
timestamp 1698431365
transform 1 0 23184 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_207
timestamp 1698431365
transform 1 0 24528 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_209
timestamp 1698431365
transform 1 0 24752 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_226
timestamp 1698431365
transform 1 0 26656 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_228
timestamp 1698431365
transform 1 0 26880 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_250
timestamp 1698431365
transform 1 0 29344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_254
timestamp 1698431365
transform 1 0 29792 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_256
timestamp 1698431365
transform 1 0 30016 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_277
timestamp 1698431365
transform 1 0 32368 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_279
timestamp 1698431365
transform 1 0 32592 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_290
timestamp 1698431365
transform 1 0 33824 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_292
timestamp 1698431365
transform 1 0 34048 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_295
timestamp 1698431365
transform 1 0 34384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_306
timestamp 1698431365
transform 1 0 35616 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_322
timestamp 1698431365
transform 1 0 37408 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_337
timestamp 1698431365
transform 1 0 39088 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_345
timestamp 1698431365
transform 1 0 39984 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_349
timestamp 1698431365
transform 1 0 40432 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_352
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_356
timestamp 1698431365
transform 1 0 41216 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_358
timestamp 1698431365
transform 1 0 41440 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_367
timestamp 1698431365
transform 1 0 42448 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_383
timestamp 1698431365
transform 1 0 44240 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_407
timestamp 1698431365
transform 1 0 46928 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_415
timestamp 1698431365
transform 1 0 47824 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_419
timestamp 1698431365
transform 1 0 48272 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_422
timestamp 1698431365
transform 1 0 48608 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_432
timestamp 1698431365
transform 1 0 49728 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_436
timestamp 1698431365
transform 1 0 50176 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_455
timestamp 1698431365
transform 1 0 52304 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_468
timestamp 1698431365
transform 1 0 53760 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_470
timestamp 1698431365
transform 1 0 53984 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_484
timestamp 1698431365
transform 1 0 55552 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_488
timestamp 1698431365
transform 1 0 56000 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_502
timestamp 1698431365
transform 1 0 57568 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_506
timestamp 1698431365
transform 1 0 58016 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_508
timestamp 1698431365
transform 1 0 58240 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_6
timestamp 1698431365
transform 1 0 2016 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_22
timestamp 1698431365
transform 1 0 3808 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_30
timestamp 1698431365
transform 1 0 4704 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_45
timestamp 1698431365
transform 1 0 6384 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_55
timestamp 1698431365
transform 1 0 7504 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_59
timestamp 1698431365
transform 1 0 7952 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_66
timestamp 1698431365
transform 1 0 8736 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_76
timestamp 1698431365
transform 1 0 9856 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_80
timestamp 1698431365
transform 1 0 10304 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_146
timestamp 1698431365
transform 1 0 17696 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_165
timestamp 1698431365
transform 1 0 19824 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_169
timestamp 1698431365
transform 1 0 20272 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_182
timestamp 1698431365
transform 1 0 21728 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_194
timestamp 1698431365
transform 1 0 23072 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_198
timestamp 1698431365
transform 1 0 23520 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_202
timestamp 1698431365
transform 1 0 23968 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_211
timestamp 1698431365
transform 1 0 24976 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_230
timestamp 1698431365
transform 1 0 27104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_234
timestamp 1698431365
transform 1 0 27552 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_238
timestamp 1698431365
transform 1 0 28000 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_242
timestamp 1698431365
transform 1 0 28448 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_249
timestamp 1698431365
transform 1 0 29232 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_281
timestamp 1698431365
transform 1 0 32816 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_285
timestamp 1698431365
transform 1 0 33264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_303
timestamp 1698431365
transform 1 0 35280 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_311
timestamp 1698431365
transform 1 0 36176 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_325
timestamp 1698431365
transform 1 0 37744 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_329
timestamp 1698431365
transform 1 0 38192 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_331
timestamp 1698431365
transform 1 0 38416 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_344
timestamp 1698431365
transform 1 0 39872 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_348
timestamp 1698431365
transform 1 0 40320 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_378
timestamp 1698431365
transform 1 0 43680 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_382
timestamp 1698431365
transform 1 0 44128 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_384
timestamp 1698431365
transform 1 0 44352 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_387
timestamp 1698431365
transform 1 0 44688 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_391
timestamp 1698431365
transform 1 0 45136 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_393
timestamp 1698431365
transform 1 0 45360 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_407
timestamp 1698431365
transform 1 0 46928 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_420
timestamp 1698431365
transform 1 0 48384 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_424
timestamp 1698431365
transform 1 0 48832 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_428
timestamp 1698431365
transform 1 0 49280 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_444
timestamp 1698431365
transform 1 0 51072 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_453
timestamp 1698431365
transform 1 0 52080 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_467
timestamp 1698431365
transform 1 0 53648 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_481
timestamp 1698431365
transform 1 0 55216 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_2
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_34
timestamp 1698431365
transform 1 0 5152 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_50
timestamp 1698431365
transform 1 0 6944 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_66
timestamp 1698431365
transform 1 0 8736 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_80
timestamp 1698431365
transform 1 0 10304 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_82
timestamp 1698431365
transform 1 0 10528 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_91
timestamp 1698431365
transform 1 0 11536 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_139
timestamp 1698431365
transform 1 0 16912 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_157
timestamp 1698431365
transform 1 0 18928 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_176
timestamp 1698431365
transform 1 0 21056 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_207
timestamp 1698431365
transform 1 0 24528 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_209
timestamp 1698431365
transform 1 0 24752 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_212
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_219
timestamp 1698431365
transform 1 0 25872 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_221
timestamp 1698431365
transform 1 0 26096 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_252
timestamp 1698431365
transform 1 0 29568 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_256
timestamp 1698431365
transform 1 0 30016 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_267
timestamp 1698431365
transform 1 0 31248 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_275
timestamp 1698431365
transform 1 0 32144 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_279
timestamp 1698431365
transform 1 0 32592 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_282
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_286
timestamp 1698431365
transform 1 0 33376 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_290
timestamp 1698431365
transform 1 0 33824 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_294
timestamp 1698431365
transform 1 0 34272 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_311
timestamp 1698431365
transform 1 0 36176 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_327
timestamp 1698431365
transform 1 0 37968 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_335
timestamp 1698431365
transform 1 0 38864 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_339
timestamp 1698431365
transform 1 0 39312 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_341
timestamp 1698431365
transform 1 0 39536 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_352
timestamp 1698431365
transform 1 0 40768 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_369
timestamp 1698431365
transform 1 0 42672 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_377
timestamp 1698431365
transform 1 0 43568 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_381
timestamp 1698431365
transform 1 0 44016 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_405
timestamp 1698431365
transform 1 0 46704 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_417
timestamp 1698431365
transform 1 0 48048 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_419
timestamp 1698431365
transform 1 0 48272 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_442
timestamp 1698431365
transform 1 0 50848 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_444
timestamp 1698431365
transform 1 0 51072 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_452
timestamp 1698431365
transform 1 0 51968 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_454
timestamp 1698431365
transform 1 0 52192 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_460
timestamp 1698431365
transform 1 0 52864 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_476
timestamp 1698431365
transform 1 0 54656 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_484
timestamp 1698431365
transform 1 0 55552 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_488
timestamp 1698431365
transform 1 0 56000 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_492
timestamp 1698431365
transform 1 0 56448 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_508
timestamp 1698431365
transform 1 0 58240 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_6
timestamp 1698431365
transform 1 0 2016 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_22
timestamp 1698431365
transform 1 0 3808 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_30
timestamp 1698431365
transform 1 0 4704 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1698431365
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_37
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_45
timestamp 1698431365
transform 1 0 6384 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_49
timestamp 1698431365
transform 1 0 6832 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_65
timestamp 1698431365
transform 1 0 8624 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_77
timestamp 1698431365
transform 1 0 9968 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_107
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_109
timestamp 1698431365
transform 1 0 13552 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_143
timestamp 1698431365
transform 1 0 17360 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_173
timestamp 1698431365
transform 1 0 20720 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_185
timestamp 1698431365
transform 1 0 22064 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_241
timestamp 1698431365
transform 1 0 28336 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_264
timestamp 1698431365
transform 1 0 30912 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_273
timestamp 1698431365
transform 1 0 31920 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_275
timestamp 1698431365
transform 1 0 32144 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_281
timestamp 1698431365
transform 1 0 32816 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_317
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_319
timestamp 1698431365
transform 1 0 37072 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_334
timestamp 1698431365
transform 1 0 38752 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_338
timestamp 1698431365
transform 1 0 39200 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_354
timestamp 1698431365
transform 1 0 40992 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_373
timestamp 1698431365
transform 1 0 43120 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_381
timestamp 1698431365
transform 1 0 44016 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_402
timestamp 1698431365
transform 1 0 46368 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_410
timestamp 1698431365
transform 1 0 47264 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_414
timestamp 1698431365
transform 1 0 47712 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_425
timestamp 1698431365
transform 1 0 48944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_427
timestamp 1698431365
transform 1 0 49168 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_454
timestamp 1698431365
transform 1 0 52192 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_469
timestamp 1698431365
transform 1 0 53872 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_477
timestamp 1698431365
transform 1 0 54768 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_481
timestamp 1698431365
transform 1 0 55216 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_2
timestamp 1698431365
transform 1 0 1568 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_34
timestamp 1698431365
transform 1 0 5152 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_42
timestamp 1698431365
transform 1 0 6048 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_62
timestamp 1698431365
transform 1 0 8288 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_92
timestamp 1698431365
transform 1 0 11648 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_94
timestamp 1698431365
transform 1 0 11872 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_124
timestamp 1698431365
transform 1 0 15232 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_138
timestamp 1698431365
transform 1 0 16800 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_187
timestamp 1698431365
transform 1 0 22288 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_207
timestamp 1698431365
transform 1 0 24528 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_209
timestamp 1698431365
transform 1 0 24752 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_227
timestamp 1698431365
transform 1 0 26768 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_231
timestamp 1698431365
transform 1 0 27216 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_250
timestamp 1698431365
transform 1 0 29344 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_257
timestamp 1698431365
transform 1 0 30128 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_261
timestamp 1698431365
transform 1 0 30576 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_265
timestamp 1698431365
transform 1 0 31024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_269
timestamp 1698431365
transform 1 0 31472 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_277
timestamp 1698431365
transform 1 0 32368 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_279
timestamp 1698431365
transform 1 0 32592 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_282
timestamp 1698431365
transform 1 0 32928 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_284
timestamp 1698431365
transform 1 0 33152 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_287
timestamp 1698431365
transform 1 0 33488 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_291
timestamp 1698431365
transform 1 0 33936 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_301
timestamp 1698431365
transform 1 0 35056 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_309
timestamp 1698431365
transform 1 0 35952 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_311
timestamp 1698431365
transform 1 0 36176 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_335
timestamp 1698431365
transform 1 0 38864 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_343
timestamp 1698431365
transform 1 0 39760 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_347
timestamp 1698431365
transform 1 0 40208 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_349
timestamp 1698431365
transform 1 0 40432 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_358
timestamp 1698431365
transform 1 0 41440 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_407
timestamp 1698431365
transform 1 0 46928 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_415
timestamp 1698431365
transform 1 0 47824 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_419
timestamp 1698431365
transform 1 0 48272 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_422
timestamp 1698431365
transform 1 0 48608 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_424
timestamp 1698431365
transform 1 0 48832 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_431
timestamp 1698431365
transform 1 0 49616 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_435
timestamp 1698431365
transform 1 0 50064 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_443
timestamp 1698431365
transform 1 0 50960 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_450
timestamp 1698431365
transform 1 0 51744 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_464
timestamp 1698431365
transform 1 0 53312 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_485
timestamp 1698431365
transform 1 0 55664 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_489
timestamp 1698431365
transform 1 0 56112 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_498
timestamp 1698431365
transform 1 0 57120 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_506
timestamp 1698431365
transform 1 0 58016 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_508
timestamp 1698431365
transform 1 0 58240 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_2
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1698431365
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_37
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_45
timestamp 1698431365
transform 1 0 6384 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_49
timestamp 1698431365
transform 1 0 6832 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_51
timestamp 1698431365
transform 1 0 7056 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_62
timestamp 1698431365
transform 1 0 8288 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_70
timestamp 1698431365
transform 1 0 9184 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_74
timestamp 1698431365
transform 1 0 9632 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_81
timestamp 1698431365
transform 1 0 10416 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_107
timestamp 1698431365
transform 1 0 13328 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_111
timestamp 1698431365
transform 1 0 13776 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_115
timestamp 1698431365
transform 1 0 14224 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_163
timestamp 1698431365
transform 1 0 19600 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_169
timestamp 1698431365
transform 1 0 20272 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_173
timestamp 1698431365
transform 1 0 20720 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_185
timestamp 1698431365
transform 1 0 22064 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_189
timestamp 1698431365
transform 1 0 22512 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_193
timestamp 1698431365
transform 1 0 22960 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_196
timestamp 1698431365
transform 1 0 23296 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_241
timestamp 1698431365
transform 1 0 28336 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_258
timestamp 1698431365
transform 1 0 30240 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_260
timestamp 1698431365
transform 1 0 30464 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_310
timestamp 1698431365
transform 1 0 36064 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_314
timestamp 1698431365
transform 1 0 36512 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_317
timestamp 1698431365
transform 1 0 36848 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_348
timestamp 1698431365
transform 1 0 40320 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_350
timestamp 1698431365
transform 1 0 40544 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_360
timestamp 1698431365
transform 1 0 41664 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_368
timestamp 1698431365
transform 1 0 42560 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_379
timestamp 1698431365
transform 1 0 43792 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_383
timestamp 1698431365
transform 1 0 44240 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_401
timestamp 1698431365
transform 1 0 46256 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_414
timestamp 1698431365
transform 1 0 47712 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_430
timestamp 1698431365
transform 1 0 49504 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_434
timestamp 1698431365
transform 1 0 49952 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_448
timestamp 1698431365
transform 1 0 51520 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_452
timestamp 1698431365
transform 1 0 51968 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_454
timestamp 1698431365
transform 1 0 52192 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_457
timestamp 1698431365
transform 1 0 52528 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_461
timestamp 1698431365
transform 1 0 52976 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_481
timestamp 1698431365
transform 1 0 55216 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_2
timestamp 1698431365
transform 1 0 1568 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_34
timestamp 1698431365
transform 1 0 5152 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_50
timestamp 1698431365
transform 1 0 6944 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_60
timestamp 1698431365
transform 1 0 8064 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_68
timestamp 1698431365
transform 1 0 8960 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_72
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_100
timestamp 1698431365
transform 1 0 12544 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_109
timestamp 1698431365
transform 1 0 13552 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_116
timestamp 1698431365
transform 1 0 14336 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_122
timestamp 1698431365
transform 1 0 15008 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_126
timestamp 1698431365
transform 1 0 15456 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_130
timestamp 1698431365
transform 1 0 15904 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_136
timestamp 1698431365
transform 1 0 16576 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_148
timestamp 1698431365
transform 1 0 17920 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_152
timestamp 1698431365
transform 1 0 18368 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_156
timestamp 1698431365
transform 1 0 18816 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_160
timestamp 1698431365
transform 1 0 19264 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_175
timestamp 1698431365
transform 1 0 20944 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_179
timestamp 1698431365
transform 1 0 21392 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_183
timestamp 1698431365
transform 1 0 21840 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_187
timestamp 1698431365
transform 1 0 22288 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_191
timestamp 1698431365
transform 1 0 22736 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_194
timestamp 1698431365
transform 1 0 23072 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_196
timestamp 1698431365
transform 1 0 23296 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_199
timestamp 1698431365
transform 1 0 23632 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_212
timestamp 1698431365
transform 1 0 25088 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_216
timestamp 1698431365
transform 1 0 25536 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_220
timestamp 1698431365
transform 1 0 25984 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_256
timestamp 1698431365
transform 1 0 30016 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_288
timestamp 1698431365
transform 1 0 33600 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_290
timestamp 1698431365
transform 1 0 33824 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_299
timestamp 1698431365
transform 1 0 34832 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_316
timestamp 1698431365
transform 1 0 36736 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_324
timestamp 1698431365
transform 1 0 37632 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_328
timestamp 1698431365
transform 1 0 38080 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_331
timestamp 1698431365
transform 1 0 38416 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_339
timestamp 1698431365
transform 1 0 39312 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_343
timestamp 1698431365
transform 1 0 39760 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_352
timestamp 1698431365
transform 1 0 40768 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_369
timestamp 1698431365
transform 1 0 42672 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_385
timestamp 1698431365
transform 1 0 44464 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_387
timestamp 1698431365
transform 1 0 44688 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_398
timestamp 1698431365
transform 1 0 45920 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_402
timestamp 1698431365
transform 1 0 46368 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_415
timestamp 1698431365
transform 1 0 47824 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_419
timestamp 1698431365
transform 1 0 48272 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_450
timestamp 1698431365
transform 1 0 51744 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_458
timestamp 1698431365
transform 1 0 52640 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_462
timestamp 1698431365
transform 1 0 53088 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_464
timestamp 1698431365
transform 1 0 53312 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_489
timestamp 1698431365
transform 1 0 56112 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_492
timestamp 1698431365
transform 1 0 56448 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_508
timestamp 1698431365
transform 1 0 58240 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_2
timestamp 1698431365
transform 1 0 1568 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_34
timestamp 1698431365
transform 1 0 5152 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_37
timestamp 1698431365
transform 1 0 5488 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_39
timestamp 1698431365
transform 1 0 5712 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_101
timestamp 1698431365
transform 1 0 12656 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_149
timestamp 1698431365
transform 1 0 18032 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_153
timestamp 1698431365
transform 1 0 18480 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_166
timestamp 1698431365
transform 1 0 19936 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_190
timestamp 1698431365
transform 1 0 22624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_192
timestamp 1698431365
transform 1 0 22848 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_195
timestamp 1698431365
transform 1 0 23184 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_219
timestamp 1698431365
transform 1 0 25872 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_221
timestamp 1698431365
transform 1 0 26096 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_241
timestamp 1698431365
transform 1 0 28336 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_252
timestamp 1698431365
transform 1 0 29568 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_262
timestamp 1698431365
transform 1 0 30688 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_264
timestamp 1698431365
transform 1 0 30912 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_288
timestamp 1698431365
transform 1 0 33600 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_292
timestamp 1698431365
transform 1 0 34048 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_296
timestamp 1698431365
transform 1 0 34496 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_306
timestamp 1698431365
transform 1 0 35616 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_314
timestamp 1698431365
transform 1 0 36512 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_317
timestamp 1698431365
transform 1 0 36848 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_325
timestamp 1698431365
transform 1 0 37744 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_329
timestamp 1698431365
transform 1 0 38192 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_331
timestamp 1698431365
transform 1 0 38416 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_340
timestamp 1698431365
transform 1 0 39424 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_348
timestamp 1698431365
transform 1 0 40320 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_352
timestamp 1698431365
transform 1 0 40768 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_354
timestamp 1698431365
transform 1 0 40992 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_361
timestamp 1698431365
transform 1 0 41776 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_377
timestamp 1698431365
transform 1 0 43568 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_402
timestamp 1698431365
transform 1 0 46368 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_418
timestamp 1698431365
transform 1 0 48160 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_425
timestamp 1698431365
transform 1 0 48944 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_429
timestamp 1698431365
transform 1 0 49392 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_433
timestamp 1698431365
transform 1 0 49840 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_449
timestamp 1698431365
transform 1 0 51632 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_453
timestamp 1698431365
transform 1 0 52080 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_457
timestamp 1698431365
transform 1 0 52528 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_489
timestamp 1698431365
transform 1 0 56112 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_505
timestamp 1698431365
transform 1 0 57904 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_55_2
timestamp 1698431365
transform 1 0 1568 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_34
timestamp 1698431365
transform 1 0 5152 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_42
timestamp 1698431365
transform 1 0 6048 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_46
timestamp 1698431365
transform 1 0 6496 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_53
timestamp 1698431365
transform 1 0 7280 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_61
timestamp 1698431365
transform 1 0 8176 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_69
timestamp 1698431365
transform 1 0 9072 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_72
timestamp 1698431365
transform 1 0 9408 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_97
timestamp 1698431365
transform 1 0 12208 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_101
timestamp 1698431365
transform 1 0 12656 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_103
timestamp 1698431365
transform 1 0 12880 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_106
timestamp 1698431365
transform 1 0 13216 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_110
timestamp 1698431365
transform 1 0 13664 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_125
timestamp 1698431365
transform 1 0 15344 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_129
timestamp 1698431365
transform 1 0 15792 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_172
timestamp 1698431365
transform 1 0 20608 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_174
timestamp 1698431365
transform 1 0 20832 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_208
timestamp 1698431365
transform 1 0 24640 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_220
timestamp 1698431365
transform 1 0 25984 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_224
timestamp 1698431365
transform 1 0 26432 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_227
timestamp 1698431365
transform 1 0 26768 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_231
timestamp 1698431365
transform 1 0 27216 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_243
timestamp 1698431365
transform 1 0 28560 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_245
timestamp 1698431365
transform 1 0 28784 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_282
timestamp 1698431365
transform 1 0 32928 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_286
timestamp 1698431365
transform 1 0 33376 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_294
timestamp 1698431365
transform 1 0 34272 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_296
timestamp 1698431365
transform 1 0 34496 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_307
timestamp 1698431365
transform 1 0 35728 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_325
timestamp 1698431365
transform 1 0 37744 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_329
timestamp 1698431365
transform 1 0 38192 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_339
timestamp 1698431365
transform 1 0 39312 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_341
timestamp 1698431365
transform 1 0 39536 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_383
timestamp 1698431365
transform 1 0 44240 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_387
timestamp 1698431365
transform 1 0 44688 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_402
timestamp 1698431365
transform 1 0 46368 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_418
timestamp 1698431365
transform 1 0 48160 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_444
timestamp 1698431365
transform 1 0 51072 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_448
timestamp 1698431365
transform 1 0 51520 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_470
timestamp 1698431365
transform 1 0 53984 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_486
timestamp 1698431365
transform 1 0 55776 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_492
timestamp 1698431365
transform 1 0 56448 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_508
timestamp 1698431365
transform 1 0 58240 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_2
timestamp 1698431365
transform 1 0 1568 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_34
timestamp 1698431365
transform 1 0 5152 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_37
timestamp 1698431365
transform 1 0 5488 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_45
timestamp 1698431365
transform 1 0 6384 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_49
timestamp 1698431365
transform 1 0 6832 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_51
timestamp 1698431365
transform 1 0 7056 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_56
timestamp 1698431365
transform 1 0 7616 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_64
timestamp 1698431365
transform 1 0 8512 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_67
timestamp 1698431365
transform 1 0 8848 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_79
timestamp 1698431365
transform 1 0 10192 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_81
timestamp 1698431365
transform 1 0 10416 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_92
timestamp 1698431365
transform 1 0 11648 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_96
timestamp 1698431365
transform 1 0 12096 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_146
timestamp 1698431365
transform 1 0 17696 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_162
timestamp 1698431365
transform 1 0 19488 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_164
timestamp 1698431365
transform 1 0 19712 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_210
timestamp 1698431365
transform 1 0 24864 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_232
timestamp 1698431365
transform 1 0 27328 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_234
timestamp 1698431365
transform 1 0 27552 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_255
timestamp 1698431365
transform 1 0 29904 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_257
timestamp 1698431365
transform 1 0 30128 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_277
timestamp 1698431365
transform 1 0 32368 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_283
timestamp 1698431365
transform 1 0 33040 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_295
timestamp 1698431365
transform 1 0 34384 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_297
timestamp 1698431365
transform 1 0 34608 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_313
timestamp 1698431365
transform 1 0 36400 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_317
timestamp 1698431365
transform 1 0 36848 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_330
timestamp 1698431365
transform 1 0 38304 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_334
timestamp 1698431365
transform 1 0 38752 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_336
timestamp 1698431365
transform 1 0 38976 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_341
timestamp 1698431365
transform 1 0 39536 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_345
timestamp 1698431365
transform 1 0 39984 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_365
timestamp 1698431365
transform 1 0 42224 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_373
timestamp 1698431365
transform 1 0 43120 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_387
timestamp 1698431365
transform 1 0 44688 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_389
timestamp 1698431365
transform 1 0 44912 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_400
timestamp 1698431365
transform 1 0 46144 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_453
timestamp 1698431365
transform 1 0 52080 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_469
timestamp 1698431365
transform 1 0 53872 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_501
timestamp 1698431365
transform 1 0 57456 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_28
timestamp 1698431365
transform 1 0 4480 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_44
timestamp 1698431365
transform 1 0 6272 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_52
timestamp 1698431365
transform 1 0 7168 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_54
timestamp 1698431365
transform 1 0 7392 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_72
timestamp 1698431365
transform 1 0 9408 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_74
timestamp 1698431365
transform 1 0 9632 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_199
timestamp 1698431365
transform 1 0 23632 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_203
timestamp 1698431365
transform 1 0 24080 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_206
timestamp 1698431365
transform 1 0 24416 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_212
timestamp 1698431365
transform 1 0 25088 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_214
timestamp 1698431365
transform 1 0 25312 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_248
timestamp 1698431365
transform 1 0 29120 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_252
timestamp 1698431365
transform 1 0 29568 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_256
timestamp 1698431365
transform 1 0 30016 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_263
timestamp 1698431365
transform 1 0 30800 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_267
timestamp 1698431365
transform 1 0 31248 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_271
timestamp 1698431365
transform 1 0 31696 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_273
timestamp 1698431365
transform 1 0 31920 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_276
timestamp 1698431365
transform 1 0 32256 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_282
timestamp 1698431365
transform 1 0 32928 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_316
timestamp 1698431365
transform 1 0 36736 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_318
timestamp 1698431365
transform 1 0 36960 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_321
timestamp 1698431365
transform 1 0 37296 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_334
timestamp 1698431365
transform 1 0 38752 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_338
timestamp 1698431365
transform 1 0 39200 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_342
timestamp 1698431365
transform 1 0 39648 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_349
timestamp 1698431365
transform 1 0 40432 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_358
timestamp 1698431365
transform 1 0 41440 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_362
timestamp 1698431365
transform 1 0 41888 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_370
timestamp 1698431365
transform 1 0 42784 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_374
timestamp 1698431365
transform 1 0 43232 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_385
timestamp 1698431365
transform 1 0 44464 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_389
timestamp 1698431365
transform 1 0 44912 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_403
timestamp 1698431365
transform 1 0 46480 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_417
timestamp 1698431365
transform 1 0 48048 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_419
timestamp 1698431365
transform 1 0 48272 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_422
timestamp 1698431365
transform 1 0 48608 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_444
timestamp 1698431365
transform 1 0 51072 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_466
timestamp 1698431365
transform 1 0 53536 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_482
timestamp 1698431365
transform 1 0 55328 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_492
timestamp 1698431365
transform 1 0 56448 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_508
timestamp 1698431365
transform 1 0 58240 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_28
timestamp 1698431365
transform 1 0 4480 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_32
timestamp 1698431365
transform 1 0 4928 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_34
timestamp 1698431365
transform 1 0 5152 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_37
timestamp 1698431365
transform 1 0 5488 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_45
timestamp 1698431365
transform 1 0 6384 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_49
timestamp 1698431365
transform 1 0 6832 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_51
timestamp 1698431365
transform 1 0 7056 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_79
timestamp 1698431365
transform 1 0 10192 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_81
timestamp 1698431365
transform 1 0 10416 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_90
timestamp 1698431365
transform 1 0 11424 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_122
timestamp 1698431365
transform 1 0 15008 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_173
timestamp 1698431365
transform 1 0 20720 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_177
timestamp 1698431365
transform 1 0 21168 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_179
timestamp 1698431365
transform 1 0 21392 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_256
timestamp 1698431365
transform 1 0 30016 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_260
timestamp 1698431365
transform 1 0 30464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_264
timestamp 1698431365
transform 1 0 30912 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_284
timestamp 1698431365
transform 1 0 33152 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_288
timestamp 1698431365
transform 1 0 33600 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_296
timestamp 1698431365
transform 1 0 34496 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_299
timestamp 1698431365
transform 1 0 34832 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_307
timestamp 1698431365
transform 1 0 35728 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_311
timestamp 1698431365
transform 1 0 36176 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_317
timestamp 1698431365
transform 1 0 36848 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_319
timestamp 1698431365
transform 1 0 37072 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_346
timestamp 1698431365
transform 1 0 40096 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_362
timestamp 1698431365
transform 1 0 41888 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_370
timestamp 1698431365
transform 1 0 42784 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_374
timestamp 1698431365
transform 1 0 43232 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_384
timestamp 1698431365
transform 1 0 44352 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_391
timestamp 1698431365
transform 1 0 45136 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_393
timestamp 1698431365
transform 1 0 45360 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_407
timestamp 1698431365
transform 1 0 46928 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_411
timestamp 1698431365
transform 1 0 47376 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_415
timestamp 1698431365
transform 1 0 47824 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_447
timestamp 1698431365
transform 1 0 51408 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_453
timestamp 1698431365
transform 1 0 52080 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_478
timestamp 1698431365
transform 1 0 54880 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_482
timestamp 1698431365
transform 1 0 55328 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_2
timestamp 1698431365
transform 1 0 1568 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_34
timestamp 1698431365
transform 1 0 5152 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_50
timestamp 1698431365
transform 1 0 6944 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_58
timestamp 1698431365
transform 1 0 7840 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_92
timestamp 1698431365
transform 1 0 11648 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_94
timestamp 1698431365
transform 1 0 11872 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_131
timestamp 1698431365
transform 1 0 16016 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_133
timestamp 1698431365
transform 1 0 16240 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_136
timestamp 1698431365
transform 1 0 16576 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_212
timestamp 1698431365
transform 1 0 25088 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_228
timestamp 1698431365
transform 1 0 26880 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_275
timestamp 1698431365
transform 1 0 32144 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_279
timestamp 1698431365
transform 1 0 32592 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_282
timestamp 1698431365
transform 1 0 32928 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_291
timestamp 1698431365
transform 1 0 33936 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_293
timestamp 1698431365
transform 1 0 34160 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_317
timestamp 1698431365
transform 1 0 36848 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_325
timestamp 1698431365
transform 1 0 37744 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_328
timestamp 1698431365
transform 1 0 38080 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_349
timestamp 1698431365
transform 1 0 40432 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_352
timestamp 1698431365
transform 1 0 40768 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_356
timestamp 1698431365
transform 1 0 41216 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_360
timestamp 1698431365
transform 1 0 41664 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_394
timestamp 1698431365
transform 1 0 45472 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_396
timestamp 1698431365
transform 1 0 45696 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_410
timestamp 1698431365
transform 1 0 47264 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_418
timestamp 1698431365
transform 1 0 48160 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_422
timestamp 1698431365
transform 1 0 48608 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_430
timestamp 1698431365
transform 1 0 49504 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_434
timestamp 1698431365
transform 1 0 49952 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_492
timestamp 1698431365
transform 1 0 56448 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_508
timestamp 1698431365
transform 1 0 58240 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_2
timestamp 1698431365
transform 1 0 1568 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_34
timestamp 1698431365
transform 1 0 5152 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_37
timestamp 1698431365
transform 1 0 5488 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_53
timestamp 1698431365
transform 1 0 7280 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_63
timestamp 1698431365
transform 1 0 8400 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_75
timestamp 1698431365
transform 1 0 9744 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_81
timestamp 1698431365
transform 1 0 10416 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_85
timestamp 1698431365
transform 1 0 10864 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_89
timestamp 1698431365
transform 1 0 11312 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_93
timestamp 1698431365
transform 1 0 11760 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_97
timestamp 1698431365
transform 1 0 12208 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_101
timestamp 1698431365
transform 1 0 12656 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_133
timestamp 1698431365
transform 1 0 16240 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_135
timestamp 1698431365
transform 1 0 16464 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_159
timestamp 1698431365
transform 1 0 19152 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_161
timestamp 1698431365
transform 1 0 19376 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_220
timestamp 1698431365
transform 1 0 25984 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_222
timestamp 1698431365
transform 1 0 26208 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_225
timestamp 1698431365
transform 1 0 26544 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_244
timestamp 1698431365
transform 1 0 28672 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_247
timestamp 1698431365
transform 1 0 29008 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_273
timestamp 1698431365
transform 1 0 31920 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_275
timestamp 1698431365
transform 1 0 32144 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_283
timestamp 1698431365
transform 1 0 33040 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_287
timestamp 1698431365
transform 1 0 33488 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_291
timestamp 1698431365
transform 1 0 33936 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_299
timestamp 1698431365
transform 1 0 34832 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_303
timestamp 1698431365
transform 1 0 35280 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_305
timestamp 1698431365
transform 1 0 35504 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_314
timestamp 1698431365
transform 1 0 36512 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_317
timestamp 1698431365
transform 1 0 36848 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_330
timestamp 1698431365
transform 1 0 38304 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_334
timestamp 1698431365
transform 1 0 38752 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_336
timestamp 1698431365
transform 1 0 38976 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_339
timestamp 1698431365
transform 1 0 39312 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_343
timestamp 1698431365
transform 1 0 39760 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_359
timestamp 1698431365
transform 1 0 41552 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_363
timestamp 1698431365
transform 1 0 42000 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_387
timestamp 1698431365
transform 1 0 44688 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_391
timestamp 1698431365
transform 1 0 45136 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_393
timestamp 1698431365
transform 1 0 45360 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_412
timestamp 1698431365
transform 1 0 47488 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_416
timestamp 1698431365
transform 1 0 47936 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_433
timestamp 1698431365
transform 1 0 49840 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_438
timestamp 1698431365
transform 1 0 50400 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_444
timestamp 1698431365
transform 1 0 51072 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_452
timestamp 1698431365
transform 1 0 51968 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_454
timestamp 1698431365
transform 1 0 52192 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_6
timestamp 1698431365
transform 1 0 2016 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_72
timestamp 1698431365
transform 1 0 9408 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_110
timestamp 1698431365
transform 1 0 13664 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_130
timestamp 1698431365
transform 1 0 15904 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_196
timestamp 1698431365
transform 1 0 23296 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_259
timestamp 1698431365
transform 1 0 30352 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_278
timestamp 1698431365
transform 1 0 32480 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_282
timestamp 1698431365
transform 1 0 32928 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_338
timestamp 1698431365
transform 1 0 39200 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_340
timestamp 1698431365
transform 1 0 39424 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_352
timestamp 1698431365
transform 1 0 40768 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_374
timestamp 1698431365
transform 1 0 43232 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_383
timestamp 1698431365
transform 1 0 44240 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_405
timestamp 1698431365
transform 1 0 46704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_409
timestamp 1698431365
transform 1 0 47152 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_418
timestamp 1698431365
transform 1 0 48160 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_441
timestamp 1698431365
transform 1 0 50736 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_473
timestamp 1698431365
transform 1 0 54320 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_481
timestamp 1698431365
transform 1 0 55216 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_489
timestamp 1698431365
transform 1 0 56112 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_492
timestamp 1698431365
transform 1 0 56448 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_508
timestamp 1698431365
transform 1 0 58240 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_2
timestamp 1698431365
transform 1 0 1568 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_34
timestamp 1698431365
transform 1 0 5152 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_37
timestamp 1698431365
transform 1 0 5488 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_53
timestamp 1698431365
transform 1 0 7280 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_57
timestamp 1698431365
transform 1 0 7728 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_92
timestamp 1698431365
transform 1 0 11648 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_102
timestamp 1698431365
transform 1 0 12768 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_104
timestamp 1698431365
transform 1 0 12992 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_107
timestamp 1698431365
transform 1 0 13328 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_109
timestamp 1698431365
transform 1 0 13552 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_148
timestamp 1698431365
transform 1 0 17920 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_150
timestamp 1698431365
transform 1 0 18144 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_163
timestamp 1698431365
transform 1 0 19600 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_167
timestamp 1698431365
transform 1 0 20048 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_177
timestamp 1698431365
transform 1 0 21168 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_191
timestamp 1698431365
transform 1 0 22736 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_195
timestamp 1698431365
transform 1 0 23184 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_198
timestamp 1698431365
transform 1 0 23520 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_255
timestamp 1698431365
transform 1 0 29904 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_257
timestamp 1698431365
transform 1 0 30128 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_283
timestamp 1698431365
transform 1 0 33040 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_309
timestamp 1698431365
transform 1 0 35952 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_313
timestamp 1698431365
transform 1 0 36400 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_334
timestamp 1698431365
transform 1 0 38752 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_338
timestamp 1698431365
transform 1 0 39200 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_362
timestamp 1698431365
transform 1 0 41888 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_370
timestamp 1698431365
transform 1 0 42784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_372
timestamp 1698431365
transform 1 0 43008 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_384
timestamp 1698431365
transform 1 0 44352 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_400
timestamp 1698431365
transform 1 0 46144 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_406
timestamp 1698431365
transform 1 0 46816 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_410
timestamp 1698431365
transform 1 0 47264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_420
timestamp 1698431365
transform 1 0 48384 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_436
timestamp 1698431365
transform 1 0 50176 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_440
timestamp 1698431365
transform 1 0 50624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_457
timestamp 1698431365
transform 1 0 52528 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_489
timestamp 1698431365
transform 1 0 56112 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_505
timestamp 1698431365
transform 1 0 57904 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_2
timestamp 1698431365
transform 1 0 1568 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_66
timestamp 1698431365
transform 1 0 8736 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_72
timestamp 1698431365
transform 1 0 9408 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_76
timestamp 1698431365
transform 1 0 9856 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_78
timestamp 1698431365
transform 1 0 10080 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_93
timestamp 1698431365
transform 1 0 11760 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_102
timestamp 1698431365
transform 1 0 12768 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_108
timestamp 1698431365
transform 1 0 13440 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_139
timestamp 1698431365
transform 1 0 16912 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_142
timestamp 1698431365
transform 1 0 17248 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_146
timestamp 1698431365
transform 1 0 17696 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_150
timestamp 1698431365
transform 1 0 18144 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_154
timestamp 1698431365
transform 1 0 18592 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_200
timestamp 1698431365
transform 1 0 23744 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_212
timestamp 1698431365
transform 1 0 25088 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_214
timestamp 1698431365
transform 1 0 25312 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_217
timestamp 1698431365
transform 1 0 25648 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_219
timestamp 1698431365
transform 1 0 25872 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_222
timestamp 1698431365
transform 1 0 26208 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_226
timestamp 1698431365
transform 1 0 26656 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_230
timestamp 1698431365
transform 1 0 27104 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_232
timestamp 1698431365
transform 1 0 27328 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_269
timestamp 1698431365
transform 1 0 31472 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_271
timestamp 1698431365
transform 1 0 31696 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_278
timestamp 1698431365
transform 1 0 32480 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_282
timestamp 1698431365
transform 1 0 32928 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_286
timestamp 1698431365
transform 1 0 33376 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_290
timestamp 1698431365
transform 1 0 33824 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_294
timestamp 1698431365
transform 1 0 34272 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_298
timestamp 1698431365
transform 1 0 34720 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_302
timestamp 1698431365
transform 1 0 35168 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_306
timestamp 1698431365
transform 1 0 35616 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_322
timestamp 1698431365
transform 1 0 37408 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_326
timestamp 1698431365
transform 1 0 37856 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_329
timestamp 1698431365
transform 1 0 38192 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_333
timestamp 1698431365
transform 1 0 38640 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_337
timestamp 1698431365
transform 1 0 39088 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_344
timestamp 1698431365
transform 1 0 39872 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_348
timestamp 1698431365
transform 1 0 40320 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_352
timestamp 1698431365
transform 1 0 40768 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_360
timestamp 1698431365
transform 1 0 41664 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_363
timestamp 1698431365
transform 1 0 42000 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_379
timestamp 1698431365
transform 1 0 43792 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_387
timestamp 1698431365
transform 1 0 44688 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_391
timestamp 1698431365
transform 1 0 45136 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_405
timestamp 1698431365
transform 1 0 46704 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_413
timestamp 1698431365
transform 1 0 47600 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_417
timestamp 1698431365
transform 1 0 48048 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_419
timestamp 1698431365
transform 1 0 48272 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_422
timestamp 1698431365
transform 1 0 48608 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_430
timestamp 1698431365
transform 1 0 49504 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_467
timestamp 1698431365
transform 1 0 53648 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_483
timestamp 1698431365
transform 1 0 55440 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_487
timestamp 1698431365
transform 1 0 55888 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_489
timestamp 1698431365
transform 1 0 56112 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_492
timestamp 1698431365
transform 1 0 56448 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_508
timestamp 1698431365
transform 1 0 58240 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_2
timestamp 1698431365
transform 1 0 1568 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_34
timestamp 1698431365
transform 1 0 5152 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_37
timestamp 1698431365
transform 1 0 5488 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_69
timestamp 1698431365
transform 1 0 9072 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_79
timestamp 1698431365
transform 1 0 10192 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_83
timestamp 1698431365
transform 1 0 10640 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_86
timestamp 1698431365
transform 1 0 10976 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_107
timestamp 1698431365
transform 1 0 13328 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_164
timestamp 1698431365
transform 1 0 19712 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_191
timestamp 1698431365
transform 1 0 22736 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_287
timestamp 1698431365
transform 1 0 33488 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_299
timestamp 1698431365
transform 1 0 34832 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_307
timestamp 1698431365
transform 1 0 35728 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_311
timestamp 1698431365
transform 1 0 36176 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_325
timestamp 1698431365
transform 1 0 37744 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_329
timestamp 1698431365
transform 1 0 38192 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_333
timestamp 1698431365
transform 1 0 38640 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_335
timestamp 1698431365
transform 1 0 38864 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_361
timestamp 1698431365
transform 1 0 41776 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_363
timestamp 1698431365
transform 1 0 42000 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_377
timestamp 1698431365
transform 1 0 43568 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_387
timestamp 1698431365
transform 1 0 44688 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_403
timestamp 1698431365
transform 1 0 46480 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_407
timestamp 1698431365
transform 1 0 46928 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_428
timestamp 1698431365
transform 1 0 49280 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_436
timestamp 1698431365
transform 1 0 50176 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_440
timestamp 1698431365
transform 1 0 50624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_447
timestamp 1698431365
transform 1 0 51408 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_457
timestamp 1698431365
transform 1 0 52528 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_471
timestamp 1698431365
transform 1 0 54096 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_479
timestamp 1698431365
transform 1 0 54992 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_2
timestamp 1698431365
transform 1 0 1568 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_66
timestamp 1698431365
transform 1 0 8736 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_72
timestamp 1698431365
transform 1 0 9408 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_90
timestamp 1698431365
transform 1 0 11424 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_96
timestamp 1698431365
transform 1 0 12096 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_100
timestamp 1698431365
transform 1 0 12544 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_104
timestamp 1698431365
transform 1 0 12992 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_128
timestamp 1698431365
transform 1 0 15680 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_142
timestamp 1698431365
transform 1 0 17248 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_144
timestamp 1698431365
transform 1 0 17472 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_192
timestamp 1698431365
transform 1 0 22848 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_194
timestamp 1698431365
transform 1 0 23072 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_225
timestamp 1698431365
transform 1 0 26544 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_227
timestamp 1698431365
transform 1 0 26768 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_279
timestamp 1698431365
transform 1 0 32592 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_345
timestamp 1698431365
transform 1 0 39984 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_349
timestamp 1698431365
transform 1 0 40432 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_382
timestamp 1698431365
transform 1 0 44128 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_386
timestamp 1698431365
transform 1 0 44576 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_396
timestamp 1698431365
transform 1 0 45696 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_400
timestamp 1698431365
transform 1 0 46144 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_482
timestamp 1698431365
transform 1 0 55328 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_492
timestamp 1698431365
transform 1 0 56448 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_508
timestamp 1698431365
transform 1 0 58240 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_28
timestamp 1698431365
transform 1 0 4480 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_32
timestamp 1698431365
transform 1 0 4928 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_34
timestamp 1698431365
transform 1 0 5152 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_37
timestamp 1698431365
transform 1 0 5488 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_69
timestamp 1698431365
transform 1 0 9072 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_85
timestamp 1698431365
transform 1 0 10864 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_93
timestamp 1698431365
transform 1 0 11760 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_97
timestamp 1698431365
transform 1 0 12208 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_101
timestamp 1698431365
transform 1 0 12656 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_107
timestamp 1698431365
transform 1 0 13328 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_127
timestamp 1698431365
transform 1 0 15568 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_137
timestamp 1698431365
transform 1 0 16688 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_139
timestamp 1698431365
transform 1 0 16912 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_160
timestamp 1698431365
transform 1 0 19264 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_177
timestamp 1698431365
transform 1 0 21168 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_179
timestamp 1698431365
transform 1 0 21392 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_231
timestamp 1698431365
transform 1 0 27216 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_233
timestamp 1698431365
transform 1 0 27440 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_244
timestamp 1698431365
transform 1 0 28672 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_247
timestamp 1698431365
transform 1 0 29008 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_273
timestamp 1698431365
transform 1 0 31920 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_287
timestamp 1698431365
transform 1 0 33488 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_297
timestamp 1698431365
transform 1 0 34608 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_301
timestamp 1698431365
transform 1 0 35056 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_317
timestamp 1698431365
transform 1 0 36848 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_331
timestamp 1698431365
transform 1 0 38416 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_335
timestamp 1698431365
transform 1 0 38864 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_339
timestamp 1698431365
transform 1 0 39312 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_343
timestamp 1698431365
transform 1 0 39760 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_362
timestamp 1698431365
transform 1 0 41888 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_383
timestamp 1698431365
transform 1 0 44240 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_405
timestamp 1698431365
transform 1 0 46704 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_409
timestamp 1698431365
transform 1 0 47152 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_412
timestamp 1698431365
transform 1 0 47488 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_442
timestamp 1698431365
transform 1 0 50848 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_463
timestamp 1698431365
transform 1 0 53200 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_495
timestamp 1698431365
transform 1 0 56784 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_503
timestamp 1698431365
transform 1 0 57680 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_507
timestamp 1698431365
transform 1 0 58128 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_2
timestamp 1698431365
transform 1 0 1568 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_36
timestamp 1698431365
transform 1 0 5376 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_41
timestamp 1698431365
transform 1 0 5936 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_47
timestamp 1698431365
transform 1 0 6608 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_59
timestamp 1698431365
transform 1 0 7952 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_63
timestamp 1698431365
transform 1 0 8400 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_70
timestamp 1698431365
transform 1 0 9184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_72
timestamp 1698431365
transform 1 0 9408 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_77
timestamp 1698431365
transform 1 0 9968 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_89
timestamp 1698431365
transform 1 0 11312 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_95
timestamp 1698431365
transform 1 0 11984 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_99
timestamp 1698431365
transform 1 0 12432 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_101
timestamp 1698431365
transform 1 0 12656 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_104
timestamp 1698431365
transform 1 0 12992 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_108
timestamp 1698431365
transform 1 0 13440 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_112
timestamp 1698431365
transform 1 0 13888 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_116
timestamp 1698431365
transform 1 0 14336 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_120
timestamp 1698431365
transform 1 0 14784 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_124
timestamp 1698431365
transform 1 0 15232 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_128
timestamp 1698431365
transform 1 0 15680 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_132
timestamp 1698431365
transform 1 0 16128 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_138
timestamp 1698431365
transform 1 0 16800 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_142
timestamp 1698431365
transform 1 0 17248 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_145
timestamp 1698431365
transform 1 0 17584 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_149
timestamp 1698431365
transform 1 0 18032 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_153
timestamp 1698431365
transform 1 0 18480 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_172
timestamp 1698431365
transform 1 0 20608 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_174
timestamp 1698431365
transform 1 0 20832 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_203
timestamp 1698431365
transform 1 0 24080 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_223
timestamp 1698431365
transform 1 0 26320 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_225
timestamp 1698431365
transform 1 0 26544 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_236
timestamp 1698431365
transform 1 0 27776 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_246
timestamp 1698431365
transform 1 0 28896 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_250
timestamp 1698431365
transform 1 0 29344 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_253
timestamp 1698431365
transform 1 0 29680 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_255
timestamp 1698431365
transform 1 0 29904 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_300
timestamp 1698431365
transform 1 0 34944 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_304
timestamp 1698431365
transform 1 0 35392 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_308
timestamp 1698431365
transform 1 0 35840 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_312
timestamp 1698431365
transform 1 0 36288 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_316
timestamp 1698431365
transform 1 0 36736 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_320
timestamp 1698431365
transform 1 0 37184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_324
timestamp 1698431365
transform 1 0 37632 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_342
timestamp 1698431365
transform 1 0 39648 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_346
timestamp 1698431365
transform 1 0 40096 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_376
timestamp 1698431365
transform 1 0 43456 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_436
timestamp 1698431365
transform 1 0 50176 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_440
timestamp 1698431365
transform 1 0 50624 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_444
timestamp 1698431365
transform 1 0 51072 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_448
timestamp 1698431365
transform 1 0 51520 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_486
timestamp 1698431365
transform 1 0 55776 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_502
timestamp 1698431365
transform 1 0 57568 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_506
timestamp 1698431365
transform 1 0 58016 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_508
timestamp 1698431365
transform 1 0 58240 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input1
timestamp 1698431365
transform -1 0 58352 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_PS_RCOSINE2_67 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 57904 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_PS_RCOSINE2_68
timestamp 1698431365
transform 1 0 57904 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_PS_RCOSINE2_69
timestamp 1698431365
transform -1 0 7952 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_PS_RCOSINE2_70
timestamp 1698431365
transform 1 0 57904 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_PS_RCOSINE2_71
timestamp 1698431365
transform 1 0 57456 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_PS_RCOSINE2_72
timestamp 1698431365
transform -1 0 6608 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_PS_RCOSINE2_73
timestamp 1698431365
transform -1 0 2016 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_PS_RCOSINE2_74
timestamp 1698431365
transform 1 0 57904 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_PS_RCOSINE2_75
timestamp 1698431365
transform -1 0 2016 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_PS_RCOSINE2_76
timestamp 1698431365
transform -1 0 11312 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_PS_RCOSINE2_77
timestamp 1698431365
transform -1 0 2016 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_PS_RCOSINE2_78
timestamp 1698431365
transform 1 0 57904 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_PS_RCOSINE2_79
timestamp 1698431365
transform 1 0 57904 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_PS_RCOSINE2_80
timestamp 1698431365
transform -1 0 2016 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_PS_RCOSINE2_81
timestamp 1698431365
transform -1 0 2688 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_PS_RCOSINE2_82
timestamp 1698431365
transform 1 0 57904 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_PS_RCOSINE2_83
timestamp 1698431365
transform 1 0 57904 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_PS_RCOSINE2_84
timestamp 1698431365
transform 1 0 57904 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_PS_RCOSINE2_85
timestamp 1698431365
transform -1 0 55328 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_PS_RCOSINE2_86
timestamp 1698431365
transform -1 0 9968 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_PS_RCOSINE2_87
timestamp 1698431365
transform -1 0 2016 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_PS_RCOSINE2_88
timestamp 1698431365
transform -1 0 9968 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_PS_RCOSINE2_89
timestamp 1698431365
transform 1 0 57904 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_PS_RCOSINE2_90
timestamp 1698431365
transform -1 0 54432 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_PS_RCOSINE2_91
timestamp 1698431365
transform 1 0 57904 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_PS_RCOSINE2_92
timestamp 1698431365
transform -1 0 55776 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_PS_RCOSINE2_93
timestamp 1698431365
transform -1 0 5824 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_PS_RCOSINE2_94
timestamp 1698431365
transform -1 0 2016 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_PS_RCOSINE2_95
timestamp 1698431365
transform 1 0 57904 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_PS_RCOSINE2_96
timestamp 1698431365
transform -1 0 11984 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_PS_RCOSINE2_97
timestamp 1698431365
transform -1 0 5936 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  OQPSK_PS_RCOSINE2_98 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 2016 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  OQPSK_PS_RCOSINE2_99
timestamp 1698431365
transform -1 0 2016 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  OQPSK_PS_RCOSINE2_100
timestamp 1698431365
transform -1 0 2464 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  OQPSK_PS_RCOSINE2_101
timestamp 1698431365
transform -1 0 2016 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  OQPSK_PS_RCOSINE2_102
timestamp 1698431365
transform 1 0 57904 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  OQPSK_PS_RCOSINE2_103
timestamp 1698431365
transform 1 0 8512 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  OQPSK_PS_RCOSINE2_104
timestamp 1698431365
transform -1 0 2464 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 55440 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698431365
transform 1 0 47264 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698431365
transform 1 0 43792 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698431365
transform 1 0 55440 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698431365
transform 1 0 55440 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698431365
transform 1 0 55440 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698431365
transform 1 0 55440 0 1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698431365
transform 1 0 55440 0 1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698431365
transform 1 0 55440 0 1 10976
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698431365
transform 1 0 55440 0 1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698431365
transform 1 0 51184 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698431365
transform 1 0 51072 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698431365
transform -1 0 43232 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698431365
transform 1 0 55440 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698431365
transform 1 0 55440 0 1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698431365
transform 1 0 55440 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698431365
transform 1 0 47264 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698431365
transform -1 0 54656 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698431365
transform 1 0 55440 0 1 53312
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698431365
transform 1 0 55440 0 1 48608
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698431365
transform 1 0 55440 0 1 50176
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output26
timestamp 1698431365
transform 1 0 55440 0 1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output27
timestamp 1698431365
transform 1 0 55440 0 1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output28
timestamp 1698431365
transform 1 0 55440 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output29
timestamp 1698431365
transform 1 0 55440 0 1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output30
timestamp 1698431365
transform -1 0 4480 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output31
timestamp 1698431365
transform -1 0 4480 0 1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output32
timestamp 1698431365
transform -1 0 4480 0 1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output33
timestamp 1698431365
transform -1 0 4480 0 -1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output34
timestamp 1698431365
transform -1 0 4480 0 -1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output35
timestamp 1698431365
transform 1 0 28896 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output36
timestamp 1698431365
transform -1 0 4480 0 -1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output37
timestamp 1698431365
transform -1 0 4480 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output38
timestamp 1698431365
transform -1 0 4480 0 -1 48608
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output39
timestamp 1698431365
transform -1 0 4480 0 1 48608
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output40
timestamp 1698431365
transform -1 0 4480 0 1 54880
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output41
timestamp 1698431365
transform -1 0 34944 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_68 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 58576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_69
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 58576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_70
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 58576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_71
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 58576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_72
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 58576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_73
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 58576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_74
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 58576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_75
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 58576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_76
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 58576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_77
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 58576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_78
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 58576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_79
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 58576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_80
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 58576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_81
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 58576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_82
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 58576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_83
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 58576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_84
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 58576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_85
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 58576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_86
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 58576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_87
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 58576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_88
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 58576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_89
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 58576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_90
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 58576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_91
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 58576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_92
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 58576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_93
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 58576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_94
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 58576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_95
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 58576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_96
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 58576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_97
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 58576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_98
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 58576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_99
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 58576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_100
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 58576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_101
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 58576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_102
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 58576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_103
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 58576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_104
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 58576 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_105
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 58576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_106
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 58576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_107
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 58576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_108
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 58576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_109
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 58576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_110
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 58576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_111
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 58576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_112
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 58576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_113
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 58576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_114
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 58576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_115
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 58576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_116
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 58576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_117
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 58576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_118
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 58576 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_119
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 58576 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_120
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 58576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_121
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 58576 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_122
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 58576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_123
timestamp 1698431365
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698431365
transform -1 0 58576 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_124
timestamp 1698431365
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698431365
transform -1 0 58576 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_125
timestamp 1698431365
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1698431365
transform -1 0 58576 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_126
timestamp 1698431365
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1698431365
transform -1 0 58576 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_127
timestamp 1698431365
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1698431365
transform -1 0 58576 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_128
timestamp 1698431365
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1698431365
transform -1 0 58576 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_129
timestamp 1698431365
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1698431365
transform -1 0 58576 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_130
timestamp 1698431365
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1698431365
transform -1 0 58576 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_131
timestamp 1698431365
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1698431365
transform -1 0 58576 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_132
timestamp 1698431365
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1698431365
transform -1 0 58576 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_133
timestamp 1698431365
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1698431365
transform -1 0 58576 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_134
timestamp 1698431365
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1698431365
transform -1 0 58576 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_135
timestamp 1698431365
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1698431365
transform -1 0 58576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_136 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_137
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_138
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_139
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_140
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_141
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_142
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_143
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_144
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_145
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_146
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_147
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_148
timestamp 1698431365
transform 1 0 50848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_149
timestamp 1698431365
transform 1 0 54656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_150
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_151
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_152
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_153
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_154
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_155
timestamp 1698431365
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_156
timestamp 1698431365
transform 1 0 56224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_157
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_158
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_159
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_160
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_161
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_162
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_163
timestamp 1698431365
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_164
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_165
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_166
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_167
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_168
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_169
timestamp 1698431365
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_170
timestamp 1698431365
transform 1 0 56224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_171
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_172
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_173
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_174
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_175
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_176
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_177
timestamp 1698431365
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_178
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_179
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_180
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_181
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_182
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_183
timestamp 1698431365
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_184
timestamp 1698431365
transform 1 0 56224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_185
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_186
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_187
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_188
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_189
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_190
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_191
timestamp 1698431365
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_192
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_193
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_194
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_195
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_196
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_197
timestamp 1698431365
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_198
timestamp 1698431365
transform 1 0 56224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_199
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_200
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_201
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_202
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_203
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_204
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_205
timestamp 1698431365
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_206
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_207
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_208
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_209
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_210
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_211
timestamp 1698431365
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_212
timestamp 1698431365
transform 1 0 56224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_213
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_214
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_215
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_216
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_217
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_218
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_219
timestamp 1698431365
transform 1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_220
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_221
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_222
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_223
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_224
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_225
timestamp 1698431365
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_226
timestamp 1698431365
transform 1 0 56224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_227
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_228
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_229
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_230
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_231
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_232
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_233
timestamp 1698431365
transform 1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_234
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_235
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_236
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_237
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_238
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_239
timestamp 1698431365
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_240
timestamp 1698431365
transform 1 0 56224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_241
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_242
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_243
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_244
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_245
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_246
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_247
timestamp 1698431365
transform 1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_248
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_249
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_250
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_251
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_252
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_253
timestamp 1698431365
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_254
timestamp 1698431365
transform 1 0 56224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_255
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_256
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_257
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_258
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_259
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_260
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_261
timestamp 1698431365
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_262
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_263
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_264
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_265
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_266
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_267
timestamp 1698431365
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_268
timestamp 1698431365
transform 1 0 56224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_269
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_270
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_271
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_272
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_273
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_274
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_275
timestamp 1698431365
transform 1 0 52304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_276
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_277
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_278
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_279
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_280
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_281
timestamp 1698431365
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_282
timestamp 1698431365
transform 1 0 56224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_283
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_284
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_285
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_286
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_287
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_288
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_289
timestamp 1698431365
transform 1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_290
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_291
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_292
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_293
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_294
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_295
timestamp 1698431365
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_296
timestamp 1698431365
transform 1 0 56224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_297
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_298
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_299
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_300
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_301
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_302
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_303
timestamp 1698431365
transform 1 0 52304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_304
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_305
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_306
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_307
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_308
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_309
timestamp 1698431365
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_310
timestamp 1698431365
transform 1 0 56224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_311
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_312
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_313
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_314
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_315
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_316
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_317
timestamp 1698431365
transform 1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_318
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_319
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_320
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_321
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_322
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_323
timestamp 1698431365
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_324
timestamp 1698431365
transform 1 0 56224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_325
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_326
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_327
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_328
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_329
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_330
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_331
timestamp 1698431365
transform 1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_332
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_333
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_334
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_335
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_336
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_337
timestamp 1698431365
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_338
timestamp 1698431365
transform 1 0 56224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_339
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_340
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_341
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_342
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_343
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_344
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_345
timestamp 1698431365
transform 1 0 52304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_346
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_347
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_348
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_349
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_350
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_351
timestamp 1698431365
transform 1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_352
timestamp 1698431365
transform 1 0 56224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_353
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_354
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_355
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_356
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_357
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_358
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_359
timestamp 1698431365
transform 1 0 52304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_360
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_361
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_362
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_363
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_364
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_365
timestamp 1698431365
transform 1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_366
timestamp 1698431365
transform 1 0 56224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_367
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_368
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_369
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_370
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_371
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_372
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_373
timestamp 1698431365
transform 1 0 52304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_374
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_375
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_376
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_377
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_378
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_379
timestamp 1698431365
transform 1 0 48384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_380
timestamp 1698431365
transform 1 0 56224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_381
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_382
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_383
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_384
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_385
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_386
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_387
timestamp 1698431365
transform 1 0 52304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_388
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_389
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_390
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_391
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_392
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_393
timestamp 1698431365
transform 1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_394
timestamp 1698431365
transform 1 0 56224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_395
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_396
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_397
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_398
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_399
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_400
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_401
timestamp 1698431365
transform 1 0 52304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_402
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_403
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_404
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_405
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_406
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_407
timestamp 1698431365
transform 1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_408
timestamp 1698431365
transform 1 0 56224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_409
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_410
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_411
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_412
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_413
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_414
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_415
timestamp 1698431365
transform 1 0 52304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_416
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_417
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_418
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_419
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_420
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_421
timestamp 1698431365
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_422
timestamp 1698431365
transform 1 0 56224 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_423
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_424
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_425
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_426
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_427
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_428
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_429
timestamp 1698431365
transform 1 0 52304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_430
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_431
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_432
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_433
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_434
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_435
timestamp 1698431365
transform 1 0 48384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_436
timestamp 1698431365
transform 1 0 56224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_437
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_438
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_439
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_440
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_441
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_442
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_443
timestamp 1698431365
transform 1 0 52304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_444
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_445
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_446
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_447
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_448
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_449
timestamp 1698431365
transform 1 0 48384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_450
timestamp 1698431365
transform 1 0 56224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_451
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_452
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_453
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_454
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_455
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_456
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_457
timestamp 1698431365
transform 1 0 52304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_458
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_459
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_460
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_461
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_462
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_463
timestamp 1698431365
transform 1 0 48384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_464
timestamp 1698431365
transform 1 0 56224 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_465
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_466
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_467
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_468
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_469
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_470
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_471
timestamp 1698431365
transform 1 0 52304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_472
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_473
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_474
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_475
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_476
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_477
timestamp 1698431365
transform 1 0 48384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_478
timestamp 1698431365
transform 1 0 56224 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_479
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_480
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_481
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_482
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_483
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_484
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_485
timestamp 1698431365
transform 1 0 52304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_486
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_487
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_488
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_489
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_490
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_491
timestamp 1698431365
transform 1 0 48384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_492
timestamp 1698431365
transform 1 0 56224 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_493
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_494
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_495
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_496
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_497
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_498
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_499
timestamp 1698431365
transform 1 0 52304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_500
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_501
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_502
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_503
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_504
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_505
timestamp 1698431365
transform 1 0 48384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_506
timestamp 1698431365
transform 1 0 56224 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_507
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_508
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_509
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_510
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_511
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_512
timestamp 1698431365
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_513
timestamp 1698431365
transform 1 0 52304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_514
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_515
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_516
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_517
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_518
timestamp 1698431365
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_519
timestamp 1698431365
transform 1 0 48384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_520
timestamp 1698431365
transform 1 0 56224 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_521
timestamp 1698431365
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_522
timestamp 1698431365
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_523
timestamp 1698431365
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_524
timestamp 1698431365
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_525
timestamp 1698431365
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_526
timestamp 1698431365
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_527
timestamp 1698431365
transform 1 0 52304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_528
timestamp 1698431365
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_529
timestamp 1698431365
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_530
timestamp 1698431365
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_531
timestamp 1698431365
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_532
timestamp 1698431365
transform 1 0 40544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_533
timestamp 1698431365
transform 1 0 48384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_534
timestamp 1698431365
transform 1 0 56224 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_535
timestamp 1698431365
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_536
timestamp 1698431365
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_537
timestamp 1698431365
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_538
timestamp 1698431365
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_539
timestamp 1698431365
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_540
timestamp 1698431365
transform 1 0 44464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_541
timestamp 1698431365
transform 1 0 52304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_542
timestamp 1698431365
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_543
timestamp 1698431365
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_544
timestamp 1698431365
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_545
timestamp 1698431365
transform 1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_546
timestamp 1698431365
transform 1 0 40544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_547
timestamp 1698431365
transform 1 0 48384 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_548
timestamp 1698431365
transform 1 0 56224 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_549
timestamp 1698431365
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_550
timestamp 1698431365
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_551
timestamp 1698431365
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_552
timestamp 1698431365
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_553
timestamp 1698431365
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_554
timestamp 1698431365
transform 1 0 44464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_555
timestamp 1698431365
transform 1 0 52304 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_556
timestamp 1698431365
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_557
timestamp 1698431365
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_558
timestamp 1698431365
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_559
timestamp 1698431365
transform 1 0 32704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_560
timestamp 1698431365
transform 1 0 40544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_561
timestamp 1698431365
transform 1 0 48384 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_562
timestamp 1698431365
transform 1 0 56224 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_563
timestamp 1698431365
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_564
timestamp 1698431365
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_565
timestamp 1698431365
transform 1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_566
timestamp 1698431365
transform 1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_567
timestamp 1698431365
transform 1 0 36624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_568
timestamp 1698431365
transform 1 0 44464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_569
timestamp 1698431365
transform 1 0 52304 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_570
timestamp 1698431365
transform 1 0 9184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_571
timestamp 1698431365
transform 1 0 17024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_572
timestamp 1698431365
transform 1 0 24864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_573
timestamp 1698431365
transform 1 0 32704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_574
timestamp 1698431365
transform 1 0 40544 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_575
timestamp 1698431365
transform 1 0 48384 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_576
timestamp 1698431365
transform 1 0 56224 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_577
timestamp 1698431365
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_578
timestamp 1698431365
transform 1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_579
timestamp 1698431365
transform 1 0 20944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_580
timestamp 1698431365
transform 1 0 28784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_581
timestamp 1698431365
transform 1 0 36624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_582
timestamp 1698431365
transform 1 0 44464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_583
timestamp 1698431365
transform 1 0 52304 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_584
timestamp 1698431365
transform 1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_585
timestamp 1698431365
transform 1 0 17024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_586
timestamp 1698431365
transform 1 0 24864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_587
timestamp 1698431365
transform 1 0 32704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_588
timestamp 1698431365
transform 1 0 40544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_589
timestamp 1698431365
transform 1 0 48384 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_590
timestamp 1698431365
transform 1 0 56224 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_591
timestamp 1698431365
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_592
timestamp 1698431365
transform 1 0 13104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_593
timestamp 1698431365
transform 1 0 20944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_594
timestamp 1698431365
transform 1 0 28784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_595
timestamp 1698431365
transform 1 0 36624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_596
timestamp 1698431365
transform 1 0 44464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_597
timestamp 1698431365
transform 1 0 52304 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_598
timestamp 1698431365
transform 1 0 9184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_599
timestamp 1698431365
transform 1 0 17024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_600
timestamp 1698431365
transform 1 0 24864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_601
timestamp 1698431365
transform 1 0 32704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_602
timestamp 1698431365
transform 1 0 40544 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_603
timestamp 1698431365
transform 1 0 48384 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_604
timestamp 1698431365
transform 1 0 56224 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_605
timestamp 1698431365
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_606
timestamp 1698431365
transform 1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_607
timestamp 1698431365
transform 1 0 20944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_608
timestamp 1698431365
transform 1 0 28784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_609
timestamp 1698431365
transform 1 0 36624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_610
timestamp 1698431365
transform 1 0 44464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_611
timestamp 1698431365
transform 1 0 52304 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_612
timestamp 1698431365
transform 1 0 5152 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_613
timestamp 1698431365
transform 1 0 8960 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_614
timestamp 1698431365
transform 1 0 12768 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_615
timestamp 1698431365
transform 1 0 16576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_616
timestamp 1698431365
transform 1 0 20384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_617
timestamp 1698431365
transform 1 0 24192 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_618
timestamp 1698431365
transform 1 0 28000 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_619
timestamp 1698431365
transform 1 0 31808 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_620
timestamp 1698431365
transform 1 0 35616 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_621
timestamp 1698431365
transform 1 0 39424 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_622
timestamp 1698431365
transform 1 0 43232 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_623
timestamp 1698431365
transform 1 0 47040 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_624
timestamp 1698431365
transform 1 0 50848 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_625
timestamp 1698431365
transform 1 0 54656 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  wire45
timestamp 1698431365
transform 1 0 19712 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  wire46
timestamp 1698431365
transform 1 0 25200 0 1 40768
box -86 -86 758 870
<< labels >>
flabel metal3 s 59200 30240 60000 30352 0 FreeSans 448 0 0 0 BitIn
port 0 nsew signal input
flabel metal3 s 0 33600 800 33712 0 FreeSans 448 0 0 0 CLK
port 1 nsew signal input
flabel metal3 s 0 30912 800 31024 0 FreeSans 448 0 0 0 EN
port 2 nsew signal input
flabel metal3 s 59200 24864 60000 24976 0 FreeSans 448 0 0 0 I[0]
port 3 nsew signal tristate
flabel metal2 s 46368 0 46480 800 0 FreeSans 448 90 0 0 I[10]
port 4 nsew signal tristate
flabel metal2 s 43680 0 43792 800 0 FreeSans 448 90 0 0 I[11]
port 5 nsew signal tristate
flabel metal2 s 42336 0 42448 800 0 FreeSans 448 90 0 0 I[12]
port 6 nsew signal tristate
flabel metal3 s 59200 23520 60000 23632 0 FreeSans 448 0 0 0 I[1]
port 7 nsew signal tristate
flabel metal3 s 59200 21504 60000 21616 0 FreeSans 448 0 0 0 I[2]
port 8 nsew signal tristate
flabel metal3 s 59200 18144 60000 18256 0 FreeSans 448 0 0 0 I[3]
port 9 nsew signal tristate
flabel metal3 s 59200 16800 60000 16912 0 FreeSans 448 0 0 0 I[4]
port 10 nsew signal tristate
flabel metal3 s 59200 15456 60000 15568 0 FreeSans 448 0 0 0 I[5]
port 11 nsew signal tristate
flabel metal3 s 59200 11424 60000 11536 0 FreeSans 448 0 0 0 I[6]
port 12 nsew signal tristate
flabel metal3 s 59200 8736 60000 8848 0 FreeSans 448 0 0 0 I[7]
port 13 nsew signal tristate
flabel metal2 s 51072 0 51184 800 0 FreeSans 448 90 0 0 I[8]
port 14 nsew signal tristate
flabel metal2 s 50400 0 50512 800 0 FreeSans 448 90 0 0 I[9]
port 15 nsew signal tristate
flabel metal2 s 40992 59200 41104 60000 0 FreeSans 448 90 0 0 Q[0]
port 16 nsew signal tristate
flabel metal3 s 59200 34944 60000 35056 0 FreeSans 448 0 0 0 Q[10]
port 17 nsew signal tristate
flabel metal3 s 59200 32928 60000 33040 0 FreeSans 448 0 0 0 Q[11]
port 18 nsew signal tristate
flabel metal3 s 59200 35616 60000 35728 0 FreeSans 448 0 0 0 Q[12]
port 19 nsew signal tristate
flabel metal2 s 45696 59200 45808 60000 0 FreeSans 448 90 0 0 Q[1]
port 20 nsew signal tristate
flabel metal2 s 52416 59200 52528 60000 0 FreeSans 448 90 0 0 Q[2]
port 21 nsew signal tristate
flabel metal3 s 59200 53088 60000 53200 0 FreeSans 448 0 0 0 Q[3]
port 22 nsew signal tristate
flabel metal3 s 59200 50400 60000 50512 0 FreeSans 448 0 0 0 Q[4]
port 23 nsew signal tristate
flabel metal3 s 59200 49728 60000 49840 0 FreeSans 448 0 0 0 Q[5]
port 24 nsew signal tristate
flabel metal3 s 59200 44352 60000 44464 0 FreeSans 448 0 0 0 Q[6]
port 25 nsew signal tristate
flabel metal3 s 59200 43008 60000 43120 0 FreeSans 448 0 0 0 Q[7]
port 26 nsew signal tristate
flabel metal3 s 59200 40320 60000 40432 0 FreeSans 448 0 0 0 Q[8]
port 27 nsew signal tristate
flabel metal3 s 59200 37632 60000 37744 0 FreeSans 448 0 0 0 Q[9]
port 28 nsew signal tristate
flabel metal3 s 0 32928 800 33040 0 FreeSans 448 0 0 0 RST
port 29 nsew signal input
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 addI[0]
port 30 nsew signal tristate
flabel metal3 s 0 28224 800 28336 0 FreeSans 448 0 0 0 addI[1]
port 31 nsew signal tristate
flabel metal3 s 0 29568 800 29680 0 FreeSans 448 0 0 0 addI[2]
port 32 nsew signal tristate
flabel metal3 s 0 28896 800 29008 0 FreeSans 448 0 0 0 addI[3]
port 33 nsew signal tristate
flabel metal3 s 0 30240 800 30352 0 FreeSans 448 0 0 0 addI[4]
port 34 nsew signal tristate
flabel metal2 s 28896 0 29008 800 0 FreeSans 448 90 0 0 addI[5]
port 35 nsew signal tristate
flabel metal3 s 0 34944 800 35056 0 FreeSans 448 0 0 0 addQ[0]
port 36 nsew signal tristate
flabel metal3 s 0 36288 800 36400 0 FreeSans 448 0 0 0 addQ[1]
port 37 nsew signal tristate
flabel metal3 s 0 47712 800 47824 0 FreeSans 448 0 0 0 addQ[2]
port 38 nsew signal tristate
flabel metal3 s 0 48384 800 48496 0 FreeSans 448 0 0 0 addQ[3]
port 39 nsew signal tristate
flabel metal3 s 0 54432 800 54544 0 FreeSans 448 0 0 0 addQ[4]
port 40 nsew signal tristate
flabel metal2 s 30912 59200 31024 60000 0 FreeSans 448 90 0 0 addQ[5]
port 41 nsew signal tristate
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 io_oeb[0]
port 42 nsew signal tristate
flabel metal3 s 59200 28224 60000 28336 0 FreeSans 448 0 0 0 io_oeb[10]
port 43 nsew signal tristate
flabel metal3 s 59200 10080 60000 10192 0 FreeSans 448 0 0 0 io_oeb[11]
port 44 nsew signal tristate
flabel metal2 s 6048 59200 6160 60000 0 FreeSans 448 90 0 0 io_oeb[12]
port 45 nsew signal tristate
flabel metal3 s 0 38976 800 39088 0 FreeSans 448 0 0 0 io_oeb[13]
port 46 nsew signal tristate
flabel metal3 s 59200 18816 60000 18928 0 FreeSans 448 0 0 0 io_oeb[14]
port 47 nsew signal tristate
flabel metal3 s 0 17472 800 17584 0 FreeSans 448 0 0 0 io_oeb[15]
port 48 nsew signal tristate
flabel metal2 s 10752 59200 10864 60000 0 FreeSans 448 90 0 0 io_oeb[16]
port 49 nsew signal tristate
flabel metal3 s 0 51072 800 51184 0 FreeSans 448 0 0 0 io_oeb[17]
port 50 nsew signal tristate
flabel metal3 s 59200 26208 60000 26320 0 FreeSans 448 0 0 0 io_oeb[18]
port 51 nsew signal tristate
flabel metal3 s 59200 25536 60000 25648 0 FreeSans 448 0 0 0 io_oeb[19]
port 52 nsew signal tristate
flabel metal3 s 0 40992 800 41104 0 FreeSans 448 0 0 0 io_oeb[1]
port 53 nsew signal tristate
flabel metal3 s 0 35616 800 35728 0 FreeSans 448 0 0 0 io_oeb[20]
port 54 nsew signal tristate
flabel metal3 s 0 31584 800 31696 0 FreeSans 448 0 0 0 io_oeb[21]
port 55 nsew signal tristate
flabel metal3 s 59200 9408 60000 9520 0 FreeSans 448 0 0 0 io_oeb[22]
port 56 nsew signal tristate
flabel metal3 s 59200 16128 60000 16240 0 FreeSans 448 0 0 0 io_oeb[23]
port 57 nsew signal tristate
flabel metal3 s 59200 22176 60000 22288 0 FreeSans 448 0 0 0 io_oeb[24]
port 58 nsew signal tristate
flabel metal2 s 54432 59200 54544 60000 0 FreeSans 448 90 0 0 io_oeb[25]
port 59 nsew signal tristate
flabel metal2 s 9408 0 9520 800 0 FreeSans 448 90 0 0 io_oeb[26]
port 60 nsew signal tristate
flabel metal3 s 0 20832 800 20944 0 FreeSans 448 0 0 0 io_oeb[27]
port 61 nsew signal tristate
flabel metal2 s 9408 59200 9520 60000 0 FreeSans 448 90 0 0 io_oeb[28]
port 62 nsew signal tristate
flabel metal3 s 59200 8064 60000 8176 0 FreeSans 448 0 0 0 io_oeb[29]
port 63 nsew signal tristate
flabel metal3 s 0 25536 800 25648 0 FreeSans 448 0 0 0 io_oeb[2]
port 64 nsew signal tristate
flabel metal2 s 52416 0 52528 800 0 FreeSans 448 90 0 0 io_oeb[30]
port 65 nsew signal tristate
flabel metal3 s 59200 19488 60000 19600 0 FreeSans 448 0 0 0 io_oeb[31]
port 66 nsew signal tristate
flabel metal2 s 55104 59200 55216 60000 0 FreeSans 448 90 0 0 io_oeb[32]
port 67 nsew signal tristate
flabel metal2 s 4704 0 4816 800 0 FreeSans 448 90 0 0 io_oeb[33]
port 68 nsew signal tristate
flabel metal3 s 0 26880 800 26992 0 FreeSans 448 0 0 0 io_oeb[34]
port 69 nsew signal tristate
flabel metal3 s 59200 12096 60000 12208 0 FreeSans 448 0 0 0 io_oeb[35]
port 70 nsew signal tristate
flabel metal2 s 11424 59200 11536 60000 0 FreeSans 448 90 0 0 io_oeb[36]
port 71 nsew signal tristate
flabel metal2 s 5376 59200 5488 60000 0 FreeSans 448 90 0 0 io_oeb[37]
port 72 nsew signal tristate
flabel metal3 s 0 42336 800 42448 0 FreeSans 448 0 0 0 io_oeb[3]
port 73 nsew signal tristate
flabel metal3 s 59200 10752 60000 10864 0 FreeSans 448 0 0 0 io_oeb[4]
port 74 nsew signal tristate
flabel metal2 s 8736 59200 8848 60000 0 FreeSans 448 90 0 0 io_oeb[5]
port 75 nsew signal tristate
flabel metal3 s 0 36960 800 37072 0 FreeSans 448 0 0 0 io_oeb[6]
port 76 nsew signal tristate
flabel metal3 s 59200 47040 60000 47152 0 FreeSans 448 0 0 0 io_oeb[7]
port 77 nsew signal tristate
flabel metal3 s 59200 13440 60000 13552 0 FreeSans 448 0 0 0 io_oeb[8]
port 78 nsew signal tristate
flabel metal2 s 7392 59200 7504 60000 0 FreeSans 448 90 0 0 io_oeb[9]
port 79 nsew signal tristate
flabel metal4 s 4448 3076 4768 56508 0 FreeSans 1280 90 0 0 vdd
port 80 nsew power bidirectional
flabel metal4 s 35168 3076 35488 56508 0 FreeSans 1280 90 0 0 vdd
port 80 nsew power bidirectional
flabel metal4 s 19808 3076 20128 56508 0 FreeSans 1280 90 0 0 vss
port 81 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 56508 0 FreeSans 1280 90 0 0 vss
port 81 nsew ground bidirectional
rlabel metal1 29960 55664 29960 55664 0 vdd
rlabel metal1 29960 56448 29960 56448 0 vss
rlabel metal2 58184 30632 58184 30632 0 BitIn
rlabel metal3 1918 33656 1918 33656 0 CLK
rlabel metal3 1302 30968 1302 30968 0 EN
rlabel metal2 57960 25256 57960 25256 0 I[0]
rlabel metal2 46424 2086 46424 2086 0 I[10]
rlabel metal2 43736 2422 43736 2422 0 I[11]
rlabel metal2 42392 2198 42392 2198 0 I[12]
rlabel metal2 57960 23800 57960 23800 0 I[1]
rlabel metal2 57960 22008 57960 22008 0 I[2]
rlabel metal2 57960 18032 57960 18032 0 I[3]
rlabel metal2 57960 16520 57960 16520 0 I[4]
rlabel metal2 57960 15120 57960 15120 0 I[5]
rlabel metal3 58618 11480 58618 11480 0 I[6]
rlabel metal3 58632 8344 58632 8344 0 I[7]
rlabel metal2 51128 2422 51128 2422 0 I[8]
rlabel metal2 50456 2198 50456 2198 0 I[9]
rlabel metal2 41048 57610 41048 57610 0 Q[0]
rlabel metal2 55384 35616 55384 35616 0 Q[10]
rlabel metal2 57960 33208 57960 33208 0 Q[11]
rlabel metal2 57736 36904 57736 36904 0 Q[12]
rlabel metal2 45752 57778 45752 57778 0 Q[1]
rlabel metal2 52472 57610 52472 57610 0 Q[2]
rlabel metal2 57288 53368 57288 53368 0 Q[3]
rlabel metal2 57848 49728 57848 49728 0 Q[4]
rlabel metal2 57960 50232 57960 50232 0 Q[5]
rlabel metal3 58618 44408 58618 44408 0 Q[6]
rlabel metal2 57960 43008 57960 43008 0 Q[7]
rlabel metal2 57960 40824 57960 40824 0 Q[8]
rlabel metal2 57960 38696 57960 38696 0 Q[9]
rlabel metal2 1736 33096 1736 33096 0 RST
rlabel metal2 33320 31528 33320 31528 0 Reg_Delay_Q.In
rlabel metal2 40488 33376 40488 33376 0 Reg_Delay_Q.Out
rlabel metal3 36792 27160 36792 27160 0 _0000_
rlabel metal2 40264 30464 40264 30464 0 _0002_
rlabel metal2 38584 29232 38584 29232 0 _0004_
rlabel metal2 39480 34384 39480 34384 0 _0005_
rlabel metal2 33096 29064 33096 29064 0 _0006_
rlabel metal2 30744 30912 30744 30912 0 _0007_
rlabel metal2 34104 32032 34104 32032 0 _0008_
rlabel metal2 9912 30576 9912 30576 0 _0009_
rlabel metal3 18984 29176 18984 29176 0 _0010_
rlabel metal2 5656 30520 5656 30520 0 _0011_
rlabel metal2 15512 30688 15512 30688 0 _0012_
rlabel metal2 21784 30576 21784 30576 0 _0013_
rlabel metal2 25368 29904 25368 29904 0 _0014_
rlabel metal3 18620 33208 18620 33208 0 _0015_
rlabel metal2 6104 34160 6104 34160 0 _0016_
rlabel metal2 21616 34328 21616 34328 0 _0017_
rlabel metal3 14392 33152 14392 33152 0 _0018_
rlabel metal2 17192 33376 17192 33376 0 _0019_
rlabel metal2 26376 33040 26376 33040 0 _0020_
rlabel metal3 43624 29400 43624 29400 0 _0021_
rlabel metal2 43568 40824 43568 40824 0 _0022_
rlabel metal2 29176 28952 29176 28952 0 _0023_
rlabel metal2 42840 25984 42840 25984 0 _0024_
rlabel metal2 44968 15512 44968 15512 0 _0025_
rlabel metal3 22792 21560 22792 21560 0 _0026_
rlabel metal2 17416 17752 17416 17752 0 _0027_
rlabel metal2 16744 20944 16744 20944 0 _0028_
rlabel metal3 24416 21560 24416 21560 0 _0029_
rlabel metal2 33544 21168 33544 21168 0 _0030_
rlabel metal3 18704 20776 18704 20776 0 _0031_
rlabel metal2 27608 19768 27608 19768 0 _0032_
rlabel metal2 16912 15624 16912 15624 0 _0033_
rlabel metal3 20496 15512 20496 15512 0 _0034_
rlabel metal2 30688 20776 30688 20776 0 _0035_
rlabel metal2 7392 18648 7392 18648 0 _0036_
rlabel metal2 28392 22344 28392 22344 0 _0037_
rlabel metal2 29624 21280 29624 21280 0 _0038_
rlabel metal3 23184 24696 23184 24696 0 _0039_
rlabel metal2 31192 21728 31192 21728 0 _0040_
rlabel metal2 31752 20608 31752 20608 0 _0041_
rlabel metal2 20104 16072 20104 16072 0 _0042_
rlabel metal2 7672 17528 7672 17528 0 _0043_
rlabel metal2 19880 16128 19880 16128 0 _0044_
rlabel metal3 22848 8456 22848 8456 0 _0045_
rlabel metal2 21784 11256 21784 11256 0 _0046_
rlabel metal3 9800 26264 9800 26264 0 _0047_
rlabel metal2 21056 19992 21056 19992 0 _0048_
rlabel metal3 17920 5880 17920 5880 0 _0049_
rlabel metal2 21560 7896 21560 7896 0 _0050_
rlabel metal2 17528 14560 17528 14560 0 _0051_
rlabel metal2 17416 13048 17416 13048 0 _0052_
rlabel metal3 18312 7448 18312 7448 0 _0053_
rlabel metal2 16296 6048 16296 6048 0 _0054_
rlabel metal2 17976 8344 17976 8344 0 _0055_
rlabel metal3 17416 7336 17416 7336 0 _0056_
rlabel metal2 24024 7784 24024 7784 0 _0057_
rlabel metal2 11256 27888 11256 27888 0 _0058_
rlabel metal2 30408 15848 30408 15848 0 _0059_
rlabel metal2 31640 21448 31640 21448 0 _0060_
rlabel metal2 37352 22064 37352 22064 0 _0061_
rlabel metal2 37688 21280 37688 21280 0 _0062_
rlabel metal2 36120 20356 36120 20356 0 _0063_
rlabel metal2 23800 18480 23800 18480 0 _0064_
rlabel metal3 20552 18312 20552 18312 0 _0065_
rlabel metal2 28840 19208 28840 19208 0 _0066_
rlabel metal3 28392 20104 28392 20104 0 _0067_
rlabel metal2 30856 20776 30856 20776 0 _0068_
rlabel metal2 14056 27552 14056 27552 0 _0069_
rlabel metal3 30744 20272 30744 20272 0 _0070_
rlabel metal2 18760 16408 18760 16408 0 _0071_
rlabel metal3 8176 16296 8176 16296 0 _0072_
rlabel metal2 16912 10584 16912 10584 0 _0073_
rlabel metal2 19208 15960 19208 15960 0 _0074_
rlabel metal2 22120 20496 22120 20496 0 _0075_
rlabel metal2 9520 19992 9520 19992 0 _0076_
rlabel metal2 10248 19600 10248 19600 0 _0077_
rlabel metal2 22848 11592 22848 11592 0 _0078_
rlabel metal2 23352 20496 23352 20496 0 _0079_
rlabel metal2 29176 26320 29176 26320 0 _0080_
rlabel metal2 33880 20776 33880 20776 0 _0081_
rlabel metal2 36232 21560 36232 21560 0 _0082_
rlabel metal2 45304 22400 45304 22400 0 _0083_
rlabel metal2 32088 20552 32088 20552 0 _0084_
rlabel metal2 35224 22120 35224 22120 0 _0085_
rlabel metal2 35784 22736 35784 22736 0 _0086_
rlabel metal3 45360 22344 45360 22344 0 _0087_
rlabel metal2 46424 22680 46424 22680 0 _0088_
rlabel metal3 47880 23016 47880 23016 0 _0089_
rlabel metal2 49784 21840 49784 21840 0 _0090_
rlabel metal2 16408 22344 16408 22344 0 _0091_
rlabel metal3 45640 22232 45640 22232 0 _0092_
rlabel metal2 46088 20888 46088 20888 0 _0093_
rlabel metal2 42840 22456 42840 22456 0 _0094_
rlabel metal2 43288 21112 43288 21112 0 _0095_
rlabel metal2 28728 15736 28728 15736 0 _0096_
rlabel metal2 20216 8008 20216 8008 0 _0097_
rlabel metal2 19768 7672 19768 7672 0 _0098_
rlabel metal2 20328 14000 20328 14000 0 _0099_
rlabel metal2 21448 9184 21448 9184 0 _0100_
rlabel metal2 15736 22848 15736 22848 0 _0101_
rlabel metal3 19096 26936 19096 26936 0 _0102_
rlabel metal2 20440 19544 20440 19544 0 _0103_
rlabel metal2 21896 15008 21896 15008 0 _0104_
rlabel metal2 16968 23800 16968 23800 0 _0105_
rlabel metal2 10416 25368 10416 25368 0 _0106_
rlabel metal2 19432 15176 19432 15176 0 _0107_
rlabel metal3 22400 26152 22400 26152 0 _0108_
rlabel metal2 20440 12992 20440 12992 0 _0109_
rlabel metal3 20776 13496 20776 13496 0 _0110_
rlabel metal4 31640 23688 31640 23688 0 _0111_
rlabel metal3 45696 20888 45696 20888 0 _0112_
rlabel metal2 26040 25368 26040 25368 0 _0113_
rlabel metal2 45864 10416 45864 10416 0 _0114_
rlabel metal2 44072 10360 44072 10360 0 _0115_
rlabel metal2 34048 25256 34048 25256 0 _0116_
rlabel metal3 37464 23128 37464 23128 0 _0117_
rlabel metal2 19432 24472 19432 24472 0 _0118_
rlabel metal2 17752 24192 17752 24192 0 _0119_
rlabel metal2 15400 25536 15400 25536 0 _0120_
rlabel metal3 15904 23016 15904 23016 0 _0121_
rlabel metal2 16520 25424 16520 25424 0 _0122_
rlabel metal3 15400 25368 15400 25368 0 _0123_
rlabel metal2 27720 25648 27720 25648 0 _0124_
rlabel metal2 17640 27104 17640 27104 0 _0125_
rlabel metal2 18424 24976 18424 24976 0 _0126_
rlabel metal2 32424 22344 32424 22344 0 _0127_
rlabel metal2 43736 18648 43736 18648 0 _0128_
rlabel metal3 29176 16856 29176 16856 0 _0129_
rlabel metal2 24248 15512 24248 15512 0 _0130_
rlabel metal2 14056 12152 14056 12152 0 _0131_
rlabel metal4 23688 14392 23688 14392 0 _0132_
rlabel metal2 24248 29232 24248 29232 0 _0133_
rlabel metal2 31864 16744 31864 16744 0 _0134_
rlabel metal2 28280 25704 28280 25704 0 _0135_
rlabel metal3 15680 3304 15680 3304 0 _0136_
rlabel metal2 29400 15680 29400 15680 0 _0137_
rlabel metal2 28952 15624 28952 15624 0 _0138_
rlabel metal2 29288 16296 29288 16296 0 _0139_
rlabel metal3 28784 15288 28784 15288 0 _0140_
rlabel metal2 12152 14504 12152 14504 0 _0141_
rlabel metal2 8344 15176 8344 15176 0 _0142_
rlabel metal2 29904 15176 29904 15176 0 _0143_
rlabel metal2 30184 15792 30184 15792 0 _0144_
rlabel metal2 30968 18144 30968 18144 0 _0145_
rlabel metal2 31080 26152 31080 26152 0 _0146_
rlabel metal2 38752 24808 38752 24808 0 _0147_
rlabel metal2 38752 22344 38752 22344 0 _0148_
rlabel metal3 40040 17416 40040 17416 0 _0149_
rlabel metal2 37464 19544 37464 19544 0 _0150_
rlabel metal3 44408 18536 44408 18536 0 _0151_
rlabel metal2 37912 20048 37912 20048 0 _0152_
rlabel metal2 31528 17976 31528 17976 0 _0153_
rlabel metal3 30072 16184 30072 16184 0 _0154_
rlabel metal3 31836 17528 31836 17528 0 _0155_
rlabel metal2 36456 19040 36456 19040 0 _0156_
rlabel metal2 9912 25536 9912 25536 0 _0157_
rlabel metal2 40040 23520 40040 23520 0 _0158_
rlabel metal2 39256 21112 39256 21112 0 _0159_
rlabel metal3 44464 20216 44464 20216 0 _0160_
rlabel metal2 46480 20104 46480 20104 0 _0161_
rlabel metal2 40712 9744 40712 9744 0 _0162_
rlabel metal3 41216 19432 41216 19432 0 _0163_
rlabel metal3 42168 20776 42168 20776 0 _0164_
rlabel metal2 41160 21000 41160 21000 0 _0165_
rlabel metal2 42168 17808 42168 17808 0 _0166_
rlabel metal2 46312 19488 46312 19488 0 _0167_
rlabel metal2 19096 17864 19096 17864 0 _0168_
rlabel metal3 47488 20776 47488 20776 0 _0169_
rlabel metal2 49560 21168 49560 21168 0 _0170_
rlabel metal2 50624 21560 50624 21560 0 _0171_
rlabel metal2 45864 20356 45864 20356 0 _0172_
rlabel metal3 49896 19096 49896 19096 0 _0173_
rlabel metal2 23520 10808 23520 10808 0 _0174_
rlabel metal2 25928 15008 25928 15008 0 _0175_
rlabel metal3 24192 15624 24192 15624 0 _0176_
rlabel metal2 23856 15288 23856 15288 0 _0177_
rlabel metal2 18984 28280 18984 28280 0 _0178_
rlabel metal3 23856 15176 23856 15176 0 _0179_
rlabel metal2 12040 7784 12040 7784 0 _0180_
rlabel metal2 18872 16576 18872 16576 0 _0181_
rlabel metal3 12264 7448 12264 7448 0 _0182_
rlabel metal2 15400 7840 15400 7840 0 _0183_
rlabel metal3 21896 23688 21896 23688 0 _0184_
rlabel metal3 20160 13608 20160 13608 0 _0185_
rlabel metal2 22792 13552 22792 13552 0 _0186_
rlabel metal2 41552 15176 41552 15176 0 _0187_
rlabel metal2 41776 21336 41776 21336 0 _0188_
rlabel metal2 25592 28672 25592 28672 0 _0189_
rlabel metal2 42616 16800 42616 16800 0 _0190_
rlabel metal2 47544 17584 47544 17584 0 _0191_
rlabel metal2 35336 14336 35336 14336 0 _0192_
rlabel metal2 35336 15260 35336 15260 0 _0193_
rlabel metal2 11144 12712 11144 12712 0 _0194_
rlabel metal3 20328 16856 20328 16856 0 _0195_
rlabel metal2 15400 11536 15400 11536 0 _0196_
rlabel metal3 15904 16184 15904 16184 0 _0197_
rlabel metal2 15232 13944 15232 13944 0 _0198_
rlabel metal2 16408 11648 16408 11648 0 _0199_
rlabel metal2 28056 27440 28056 27440 0 _0200_
rlabel metal2 13384 15148 13384 15148 0 _0201_
rlabel metal2 8120 15792 8120 15792 0 _0202_
rlabel metal2 19880 11200 19880 11200 0 _0203_
rlabel metal2 18424 10080 18424 10080 0 _0204_
rlabel metal3 12544 10584 12544 10584 0 _0205_
rlabel metal3 14896 15288 14896 15288 0 _0206_
rlabel metal2 16632 13552 16632 13552 0 _0207_
rlabel metal3 15400 13160 15400 13160 0 _0208_
rlabel metal3 22904 1624 22904 1624 0 _0209_
rlabel metal2 35000 14224 35000 14224 0 _0210_
rlabel metal3 29344 25480 29344 25480 0 _0211_
rlabel metal2 34496 17080 34496 17080 0 _0212_
rlabel metal2 34664 15736 34664 15736 0 _0213_
rlabel metal2 33040 22904 33040 22904 0 _0214_
rlabel metal2 31752 15624 31752 15624 0 _0215_
rlabel metal3 33936 16072 33936 16072 0 _0216_
rlabel metal2 45752 16520 45752 16520 0 _0217_
rlabel metal2 20664 17192 20664 17192 0 _0218_
rlabel metal2 21224 17192 21224 17192 0 _0219_
rlabel metal2 24808 17416 24808 17416 0 _0220_
rlabel metal2 18256 25816 18256 25816 0 _0221_
rlabel metal2 31304 26096 31304 26096 0 _0222_
rlabel metal2 23464 18816 23464 18816 0 _0223_
rlabel metal2 26040 17976 26040 17976 0 _0224_
rlabel metal2 34776 17808 34776 17808 0 _0225_
rlabel metal2 39480 18368 39480 18368 0 _0226_
rlabel metal2 38472 19152 38472 19152 0 _0227_
rlabel metal2 45976 18032 45976 18032 0 _0228_
rlabel metal3 46816 17640 46816 17640 0 _0229_
rlabel metal3 48944 17640 48944 17640 0 _0230_
rlabel metal3 50400 17528 50400 17528 0 _0231_
rlabel metal3 44688 8344 44688 8344 0 _0232_
rlabel metal2 31864 25368 31864 25368 0 _0233_
rlabel metal2 43400 25424 43400 25424 0 _0234_
rlabel metal2 43736 20188 43736 20188 0 _0235_
rlabel metal2 43568 18648 43568 18648 0 _0236_
rlabel metal2 44240 19432 44240 19432 0 _0237_
rlabel metal3 44856 20440 44856 20440 0 _0238_
rlabel metal2 48888 20720 48888 20720 0 _0239_
rlabel metal2 50344 20412 50344 20412 0 _0240_
rlabel metal2 52416 19096 52416 19096 0 _0241_
rlabel metal2 47376 18200 47376 18200 0 _0242_
rlabel metal3 34160 25592 34160 25592 0 _0243_
rlabel metal2 47656 16016 47656 16016 0 _0244_
rlabel metal2 18984 12656 18984 12656 0 _0245_
rlabel metal2 17976 11536 17976 11536 0 _0246_
rlabel metal2 19544 11312 19544 11312 0 _0247_
rlabel metal2 19432 9184 19432 9184 0 _0248_
rlabel metal2 17528 8456 17528 8456 0 _0249_
rlabel metal3 16576 8232 16576 8232 0 _0250_
rlabel metal2 19656 11144 19656 11144 0 _0251_
rlabel metal2 41720 11816 41720 11816 0 _0252_
rlabel metal2 42112 13160 42112 13160 0 _0253_
rlabel metal3 36624 25256 36624 25256 0 _0254_
rlabel metal3 42336 12936 42336 12936 0 _0255_
rlabel metal2 46200 13944 46200 13944 0 _0256_
rlabel metal2 16464 9240 16464 9240 0 _0257_
rlabel metal2 30072 12544 30072 12544 0 _0258_
rlabel metal2 25256 14672 25256 14672 0 _0259_
rlabel metal3 20216 14112 20216 14112 0 _0260_
rlabel metal2 24808 14112 24808 14112 0 _0261_
rlabel metal2 21336 14056 21336 14056 0 _0262_
rlabel metal2 29400 13664 29400 13664 0 _0263_
rlabel metal3 32368 13832 32368 13832 0 _0264_
rlabel metal2 37352 25872 37352 25872 0 _0265_
rlabel metal2 41496 14168 41496 14168 0 _0266_
rlabel metal2 33432 15232 33432 15232 0 _0267_
rlabel metal2 32424 13832 32424 13832 0 _0268_
rlabel metal3 32144 15288 32144 15288 0 _0269_
rlabel metal2 41160 14616 41160 14616 0 _0270_
rlabel metal2 45024 13944 45024 13944 0 _0271_
rlabel metal2 29848 17136 29848 17136 0 _0272_
rlabel metal2 27160 18592 27160 18592 0 _0273_
rlabel metal2 29568 17640 29568 17640 0 _0274_
rlabel metal2 29960 17920 29960 17920 0 _0275_
rlabel metal2 29736 17584 29736 17584 0 _0276_
rlabel metal2 23688 14336 23688 14336 0 _0277_
rlabel metal2 34552 17696 34552 17696 0 _0278_
rlabel metal3 36792 15288 36792 15288 0 _0279_
rlabel metal2 41160 15120 41160 15120 0 _0280_
rlabel metal2 37408 18312 37408 18312 0 _0281_
rlabel metal3 17360 13720 17360 13720 0 _0282_
rlabel metal3 25200 7448 25200 7448 0 _0283_
rlabel metal2 24584 7672 24584 7672 0 _0284_
rlabel metal2 20776 10304 20776 10304 0 _0285_
rlabel metal3 8120 43512 8120 43512 0 _0286_
rlabel metal3 19656 4536 19656 4536 0 _0287_
rlabel metal2 23800 5208 23800 5208 0 _0288_
rlabel metal2 25424 13720 25424 13720 0 _0289_
rlabel metal2 24920 6888 24920 6888 0 _0290_
rlabel metal2 26488 6552 26488 6552 0 _0291_
rlabel metal2 17864 5488 17864 5488 0 _0292_
rlabel metal2 18032 5096 18032 5096 0 _0293_
rlabel metal3 24864 4424 24864 4424 0 _0294_
rlabel metal2 15288 5320 15288 5320 0 _0295_
rlabel metal2 14280 6384 14280 6384 0 _0296_
rlabel metal2 7560 43176 7560 43176 0 _0297_
rlabel metal2 13832 6216 13832 6216 0 _0298_
rlabel metal2 15176 6216 15176 6216 0 _0299_
rlabel metal2 28392 6664 28392 6664 0 _0300_
rlabel metal2 38976 13720 38976 13720 0 _0301_
rlabel metal2 44856 14056 44856 14056 0 _0302_
rlabel metal3 46312 13944 46312 13944 0 _0303_
rlabel metal2 43288 14336 43288 14336 0 _0304_
rlabel metal2 37968 15288 37968 15288 0 _0305_
rlabel metal2 43176 14560 43176 14560 0 _0306_
rlabel metal2 46200 14952 46200 14952 0 _0307_
rlabel metal2 13832 52304 13832 52304 0 _0308_
rlabel metal2 47712 13944 47712 13944 0 _0309_
rlabel metal2 50120 16016 50120 16016 0 _0310_
rlabel metal2 49560 19824 49560 19824 0 _0311_
rlabel metal2 48776 18088 48776 18088 0 _0312_
rlabel metal2 51688 17192 51688 17192 0 _0313_
rlabel metal2 51240 16800 51240 16800 0 _0314_
rlabel metal3 52136 15960 52136 15960 0 _0315_
rlabel metal2 46760 14616 46760 14616 0 _0316_
rlabel metal2 45976 14000 45976 14000 0 _0317_
rlabel metal2 8344 52808 8344 52808 0 _0318_
rlabel metal3 47936 13048 47936 13048 0 _0319_
rlabel metal2 25480 5040 25480 5040 0 _0320_
rlabel metal2 26040 4648 26040 4648 0 _0321_
rlabel metal2 25760 5208 25760 5208 0 _0322_
rlabel metal2 24472 12376 24472 12376 0 _0323_
rlabel metal2 22344 5712 22344 5712 0 _0324_
rlabel metal2 21560 5936 21560 5936 0 _0325_
rlabel metal2 26320 5880 26320 5880 0 _0326_
rlabel metal2 27048 5824 27048 5824 0 _0327_
rlabel metal2 41720 10416 41720 10416 0 _0328_
rlabel metal3 13440 52920 13440 52920 0 _0329_
rlabel metal3 42616 11368 42616 11368 0 _0330_
rlabel metal2 43848 11620 43848 11620 0 _0331_
rlabel metal2 46648 12096 46648 12096 0 _0332_
rlabel metal2 39704 14896 39704 14896 0 _0333_
rlabel metal2 27272 13104 27272 13104 0 _0334_
rlabel metal2 26376 12992 26376 12992 0 _0335_
rlabel metal2 21112 10864 21112 10864 0 _0336_
rlabel metal3 22568 10584 22568 10584 0 _0337_
rlabel metal2 27160 12264 27160 12264 0 _0338_
rlabel metal2 27048 14840 27048 14840 0 _0339_
rlabel metal3 13552 36680 13552 36680 0 _0340_
rlabel metal2 39816 14840 39816 14840 0 _0341_
rlabel metal2 36120 17528 36120 17528 0 _0342_
rlabel metal2 36008 16240 36008 16240 0 _0343_
rlabel metal3 35448 16856 35448 16856 0 _0344_
rlabel metal2 37968 16744 37968 16744 0 _0345_
rlabel metal2 39032 15568 39032 15568 0 _0346_
rlabel metal2 45640 14392 45640 14392 0 _0347_
rlabel metal2 40152 15400 40152 15400 0 _0348_
rlabel metal3 39088 15848 39088 15848 0 _0349_
rlabel metal2 39704 12208 39704 12208 0 _0350_
rlabel metal2 12264 47152 12264 47152 0 _0351_
rlabel metal2 40824 15792 40824 15792 0 _0352_
rlabel metal2 45416 15848 45416 15848 0 _0353_
rlabel metal2 46760 12432 46760 12432 0 _0354_
rlabel metal2 49224 12600 49224 12600 0 _0355_
rlabel metal2 51800 15120 51800 15120 0 _0356_
rlabel metal2 47096 15512 47096 15512 0 _0357_
rlabel metal3 45360 14280 45360 14280 0 _0358_
rlabel metal2 45920 14616 45920 14616 0 _0359_
rlabel metal3 49728 15400 49728 15400 0 _0360_
rlabel metal2 7112 40880 7112 40880 0 _0361_
rlabel metal2 51016 15624 51016 15624 0 _0362_
rlabel metal2 51352 15232 51352 15232 0 _0363_
rlabel metal2 52864 15288 52864 15288 0 _0364_
rlabel metal2 46984 11424 46984 11424 0 _0365_
rlabel metal2 49000 10864 49000 10864 0 _0366_
rlabel metal2 42392 10864 42392 10864 0 _0367_
rlabel metal3 24696 10808 24696 10808 0 _0368_
rlabel metal2 15736 6104 15736 6104 0 _0369_
rlabel metal2 23184 24696 23184 24696 0 _0370_
rlabel metal2 9016 40712 9016 40712 0 _0371_
rlabel metal3 23576 24584 23576 24584 0 _0372_
rlabel metal2 24528 10808 24528 10808 0 _0373_
rlabel metal2 28280 9520 28280 9520 0 _0374_
rlabel metal3 28672 9240 28672 9240 0 _0375_
rlabel metal2 26488 10080 26488 10080 0 _0376_
rlabel metal2 42168 10752 42168 10752 0 _0377_
rlabel metal2 47208 10192 47208 10192 0 _0378_
rlabel metal3 31920 8232 31920 8232 0 _0379_
rlabel metal3 34384 8008 34384 8008 0 _0380_
rlabel metal2 22904 4816 22904 4816 0 _0381_
rlabel metal2 13384 44072 13384 44072 0 _0382_
rlabel metal2 26600 8008 26600 8008 0 _0383_
rlabel metal2 19768 4984 19768 4984 0 _0384_
rlabel metal2 19544 4928 19544 4928 0 _0385_
rlabel metal2 19096 4648 19096 4648 0 _0386_
rlabel metal3 20720 4536 20720 4536 0 _0387_
rlabel metal2 21784 6048 21784 6048 0 _0388_
rlabel metal2 31640 9296 31640 9296 0 _0389_
rlabel metal2 44296 9184 44296 9184 0 _0390_
rlabel metal2 20440 6216 20440 6216 0 _0391_
rlabel metal2 20216 6720 20216 6720 0 _0392_
rlabel metal3 21168 49000 21168 49000 0 _0393_
rlabel metal2 22456 5824 22456 5824 0 _0394_
rlabel metal3 20440 5096 20440 5096 0 _0395_
rlabel metal2 22008 4872 22008 4872 0 _0396_
rlabel metal3 22512 19096 22512 19096 0 _0397_
rlabel metal2 22736 5096 22736 5096 0 _0398_
rlabel metal2 38248 8792 38248 8792 0 _0399_
rlabel metal2 38976 9800 38976 9800 0 _0400_
rlabel metal2 43848 9296 43848 9296 0 _0401_
rlabel metal2 45416 9744 45416 9744 0 _0402_
rlabel metal3 44632 9800 44632 9800 0 _0403_
rlabel metal2 21896 47096 21896 47096 0 _0404_
rlabel metal3 46704 9912 46704 9912 0 _0405_
rlabel metal3 48272 10584 48272 10584 0 _0406_
rlabel metal2 50792 9072 50792 9072 0 _0407_
rlabel metal2 50344 15232 50344 15232 0 _0408_
rlabel metal2 49560 13440 49560 13440 0 _0409_
rlabel metal2 50792 12376 50792 12376 0 _0410_
rlabel metal2 51352 13832 51352 13832 0 _0411_
rlabel metal2 50232 11536 50232 11536 0 _0412_
rlabel metal2 51184 11256 51184 11256 0 _0413_
rlabel metal2 11144 36680 11144 36680 0 _0414_
rlabel metal2 49336 7924 49336 7924 0 _0415_
rlabel metal2 41496 7280 41496 7280 0 _0416_
rlabel metal2 15288 6216 15288 6216 0 _0417_
rlabel metal2 18200 7560 18200 7560 0 _0418_
rlabel metal3 21896 2632 21896 2632 0 _0419_
rlabel metal3 25368 7336 25368 7336 0 _0420_
rlabel metal2 31976 7448 31976 7448 0 _0421_
rlabel metal2 42728 7952 42728 7952 0 _0422_
rlabel metal3 34608 15512 34608 15512 0 _0423_
rlabel metal2 15288 10752 15288 10752 0 _0424_
rlabel metal2 18648 34832 18648 34832 0 _0425_
rlabel metal2 15960 9072 15960 9072 0 _0426_
rlabel metal3 16408 9240 16408 9240 0 _0427_
rlabel metal2 11928 14448 11928 14448 0 _0428_
rlabel metal2 16072 12432 16072 12432 0 _0429_
rlabel metal4 18424 10864 18424 10864 0 _0430_
rlabel metal2 33320 11648 33320 11648 0 _0431_
rlabel metal2 40600 10640 40600 10640 0 _0432_
rlabel metal2 42616 9408 42616 9408 0 _0433_
rlabel metal3 44128 8232 44128 8232 0 _0434_
rlabel metal4 43736 8232 43736 8232 0 _0435_
rlabel metal3 9240 49784 9240 49784 0 _0436_
rlabel metal2 45864 8232 45864 8232 0 _0437_
rlabel metal2 35336 9296 35336 9296 0 _0438_
rlabel metal2 26040 9632 26040 9632 0 _0439_
rlabel metal2 27552 25368 27552 25368 0 _0440_
rlabel metal2 18536 9464 18536 9464 0 _0441_
rlabel metal3 21784 9016 21784 9016 0 _0442_
rlabel metal3 25256 9016 25256 9016 0 _0443_
rlabel metal2 25816 8736 25816 8736 0 _0444_
rlabel metal2 45528 7672 45528 7672 0 _0445_
rlabel metal2 48328 7056 48328 7056 0 _0446_
rlabel via2 10360 52136 10360 52136 0 _0447_
rlabel metal2 50904 7840 50904 7840 0 _0448_
rlabel metal2 50008 9296 50008 9296 0 _0449_
rlabel metal2 51072 8792 51072 8792 0 _0450_
rlabel metal2 51240 7924 51240 7924 0 _0451_
rlabel metal2 51352 7840 51352 7840 0 _0452_
rlabel metal3 46424 5880 46424 5880 0 _0453_
rlabel metal3 23464 11368 23464 11368 0 _0454_
rlabel metal2 23632 11592 23632 11592 0 _0455_
rlabel metal2 24360 11592 24360 11592 0 _0456_
rlabel metal2 11928 53480 11928 53480 0 _0457_
rlabel metal3 27384 11088 27384 11088 0 _0458_
rlabel metal2 33432 10080 33432 10080 0 _0459_
rlabel metal2 39704 10976 39704 10976 0 _0460_
rlabel metal2 33656 6888 33656 6888 0 _0461_
rlabel metal2 25144 5152 25144 5152 0 _0462_
rlabel metal2 28952 4928 28952 4928 0 _0463_
rlabel metal2 28952 4088 28952 4088 0 _0464_
rlabel metal2 26936 5376 26936 5376 0 _0465_
rlabel metal2 31640 5600 31640 5600 0 _0466_
rlabel metal2 31528 6216 31528 6216 0 _0467_
rlabel metal2 8736 52248 8736 52248 0 _0468_
rlabel metal2 31864 5432 31864 5432 0 _0469_
rlabel metal2 33432 4648 33432 4648 0 _0470_
rlabel metal2 31864 3920 31864 3920 0 _0471_
rlabel metal2 41496 10976 41496 10976 0 _0472_
rlabel metal2 23128 9800 23128 9800 0 _0473_
rlabel metal3 30688 10472 30688 10472 0 _0474_
rlabel metal2 30856 7448 30856 7448 0 _0475_
rlabel metal2 46424 5656 46424 5656 0 _0476_
rlabel metal2 48888 5936 48888 5936 0 _0477_
rlabel metal3 48720 8904 48720 8904 0 _0478_
rlabel metal2 10360 43064 10360 43064 0 _0479_
rlabel metal2 49000 7952 49000 7952 0 _0480_
rlabel metal2 48720 5992 48720 5992 0 _0481_
rlabel metal2 50512 5880 50512 5880 0 _0482_
rlabel metal3 31752 4536 31752 4536 0 _0483_
rlabel metal2 45192 5432 45192 5432 0 _0484_
rlabel metal2 47432 4480 47432 4480 0 _0485_
rlabel metal2 24696 29904 24696 29904 0 _0486_
rlabel metal3 30240 12152 30240 12152 0 _0487_
rlabel metal3 33544 11928 33544 11928 0 _0488_
rlabel metal2 10472 45472 10472 45472 0 _0489_
rlabel metal2 35056 4312 35056 4312 0 _0490_
rlabel metal2 18200 28840 18200 28840 0 _0491_
rlabel metal3 22848 26376 22848 26376 0 _0492_
rlabel metal2 27216 21112 27216 21112 0 _0493_
rlabel metal2 34776 11424 34776 11424 0 _0494_
rlabel metal2 34664 10696 34664 10696 0 _0495_
rlabel metal2 34776 10864 34776 10864 0 _0496_
rlabel metal2 34720 5096 34720 5096 0 _0497_
rlabel metal3 29904 8008 29904 8008 0 _0498_
rlabel metal2 28112 8344 28112 8344 0 _0499_
rlabel metal3 17416 37464 17416 37464 0 _0500_
rlabel metal3 29232 8120 29232 8120 0 _0501_
rlabel metal3 31752 8120 31752 8120 0 _0502_
rlabel metal2 33488 8008 33488 8008 0 _0503_
rlabel metal2 34720 5320 34720 5320 0 _0504_
rlabel metal2 35112 4704 35112 4704 0 _0505_
rlabel metal3 35000 4984 35000 4984 0 _0506_
rlabel metal2 35336 4536 35336 4536 0 _0507_
rlabel metal2 47208 4032 47208 4032 0 _0508_
rlabel metal2 50120 5376 50120 5376 0 _0509_
rlabel metal3 50176 4984 50176 4984 0 _0510_
rlabel metal2 24696 36848 24696 36848 0 _0511_
rlabel metal2 50848 4424 50848 4424 0 _0512_
rlabel metal2 50568 4536 50568 4536 0 _0513_
rlabel metal2 27496 9856 27496 9856 0 _0514_
rlabel metal2 38696 9408 38696 9408 0 _0515_
rlabel metal3 41272 8008 41272 8008 0 _0516_
rlabel metal2 39536 9016 39536 9016 0 _0517_
rlabel metal2 39144 5992 39144 5992 0 _0518_
rlabel metal2 32648 6720 32648 6720 0 _0519_
rlabel metal2 35336 7392 35336 7392 0 _0520_
rlabel metal3 25144 56168 25144 56168 0 _0521_
rlabel metal2 35896 6440 35896 6440 0 _0522_
rlabel metal2 38472 4816 38472 4816 0 _0523_
rlabel metal2 35896 12320 35896 12320 0 _0524_
rlabel metal2 36960 6664 36960 6664 0 _0525_
rlabel via2 39032 5096 39032 5096 0 _0526_
rlabel metal2 38808 4648 38808 4648 0 _0527_
rlabel metal3 36288 4200 36288 4200 0 _0528_
rlabel metal3 44800 4872 44800 4872 0 _0529_
rlabel metal2 46536 5376 46536 5376 0 _0530_
rlabel metal2 49336 5096 49336 5096 0 _0531_
rlabel metal2 14952 54880 14952 54880 0 _0532_
rlabel metal3 47432 5208 47432 5208 0 _0533_
rlabel metal2 46200 5320 46200 5320 0 _0534_
rlabel metal3 46592 5096 46592 5096 0 _0535_
rlabel metal2 40040 5824 40040 5824 0 _0536_
rlabel metal2 40600 5432 40600 5432 0 _0537_
rlabel metal2 24248 9744 24248 9744 0 _0538_
rlabel metal2 24136 9912 24136 9912 0 _0539_
rlabel metal2 24472 9968 24472 9968 0 _0540_
rlabel metal2 36344 11088 36344 11088 0 _0541_
rlabel metal2 19152 45864 19152 45864 0 _0542_
rlabel metal2 37912 11424 37912 11424 0 _0543_
rlabel metal2 37688 10696 37688 10696 0 _0544_
rlabel metal2 38864 6664 38864 6664 0 _0545_
rlabel metal2 39480 5432 39480 5432 0 _0546_
rlabel metal2 41496 6104 41496 6104 0 _0547_
rlabel metal2 41328 5096 41328 5096 0 _0548_
rlabel metal2 43064 5040 43064 5040 0 _0549_
rlabel metal2 42952 4928 42952 4928 0 _0550_
rlabel metal2 42168 5544 42168 5544 0 _0551_
rlabel metal2 43288 5488 43288 5488 0 _0552_
rlabel metal3 25144 40264 25144 40264 0 _0553_
rlabel metal2 43400 4648 43400 4648 0 _0554_
rlabel metal2 39144 7056 39144 7056 0 _0555_
rlabel metal2 38584 7448 38584 7448 0 _0556_
rlabel metal2 39032 7728 39032 7728 0 _0557_
rlabel metal2 44184 5600 44184 5600 0 _0558_
rlabel metal2 42840 6776 42840 6776 0 _0559_
rlabel metal2 40040 5208 40040 5208 0 _0560_
rlabel metal2 42224 6104 42224 6104 0 _0561_
rlabel metal3 25704 36176 25704 36176 0 _0562_
rlabel metal2 49784 23464 49784 23464 0 _0563_
rlabel metal2 33544 29288 33544 29288 0 _0564_
rlabel metal2 31416 30072 31416 30072 0 _0565_
rlabel metal3 26712 9240 26712 9240 0 _0566_
rlabel metal2 25816 31360 25816 31360 0 _0567_
rlabel metal2 33768 31248 33768 31248 0 _0568_
rlabel metal2 23184 55944 23184 55944 0 _0569_
rlabel metal2 17864 31024 17864 31024 0 _0570_
rlabel metal2 10136 29680 10136 29680 0 _0571_
rlabel metal3 20552 34104 20552 34104 0 _0572_
rlabel metal2 18312 29400 18312 29400 0 _0573_
rlabel metal3 20272 29288 20272 29288 0 _0574_
rlabel metal3 16044 30072 16044 30072 0 _0575_
rlabel metal3 21056 29512 21056 29512 0 _0576_
rlabel metal2 20160 51352 20160 51352 0 _0577_
rlabel metal3 16576 30184 16576 30184 0 _0578_
rlabel metal2 22232 29176 22232 29176 0 _0579_
rlabel metal2 21448 29344 21448 29344 0 _0580_
rlabel metal2 24024 29960 24024 29960 0 _0581_
rlabel metal3 19208 32648 19208 32648 0 _0582_
rlabel metal3 23912 32312 23912 32312 0 _0583_
rlabel metal2 25704 29680 25704 29680 0 _0584_
rlabel metal3 33544 39032 33544 39032 0 _0585_
rlabel metal2 19936 33320 19936 33320 0 _0586_
rlabel metal3 23856 33320 23856 33320 0 _0587_
rlabel metal2 22792 33040 22792 33040 0 _0588_
rlabel metal2 25592 32816 25592 32816 0 _0589_
rlabel metal2 26376 33992 26376 33992 0 _0590_
rlabel metal2 25256 33600 25256 33600 0 _0591_
rlabel metal2 14504 54152 14504 54152 0 _0592_
rlabel metal2 26488 33656 26488 33656 0 _0593_
rlabel metal3 44968 30072 44968 30072 0 _0594_
rlabel metal2 31808 28616 31808 28616 0 _0595_
rlabel metal3 30296 28616 30296 28616 0 _0596_
rlabel metal2 43064 25368 43064 25368 0 _0597_
rlabel metal3 14616 55216 14616 55216 0 _0598_
rlabel metal2 10472 51296 10472 51296 0 _0599_
rlabel metal2 7672 46144 7672 46144 0 _0600_
rlabel metal2 18760 46536 18760 46536 0 _0601_
rlabel metal2 19432 46648 19432 46648 0 _0602_
rlabel metal3 33096 46872 33096 46872 0 _0603_
rlabel metal3 34328 45528 34328 45528 0 _0604_
rlabel metal2 39816 37352 39816 37352 0 _0605_
rlabel metal2 35112 21056 35112 21056 0 _0606_
rlabel metal2 36568 19208 36568 19208 0 _0607_
rlabel metal2 37184 26824 37184 26824 0 _0608_
rlabel metal2 22008 28672 22008 28672 0 _0609_
rlabel metal3 41160 24584 41160 24584 0 _0610_
rlabel metal2 37464 24584 37464 24584 0 _0611_
rlabel metal2 38696 28112 38696 28112 0 _0612_
rlabel metal2 38192 27608 38192 27608 0 _0613_
rlabel metal2 35672 28280 35672 28280 0 _0614_
rlabel metal2 37464 27272 37464 27272 0 _0615_
rlabel metal2 39424 53256 39424 53256 0 _0616_
rlabel metal2 39088 45752 39088 45752 0 _0617_
rlabel metal2 41832 39144 41832 39144 0 _0618_
rlabel metal2 38696 31836 38696 31836 0 _0619_
rlabel metal3 40376 31192 40376 31192 0 _0620_
rlabel metal2 39088 30744 39088 30744 0 _0621_
rlabel metal3 40600 30968 40600 30968 0 _0622_
rlabel metal2 39480 29512 39480 29512 0 _0623_
rlabel metal2 34496 49224 34496 49224 0 _0624_
rlabel metal2 9184 50568 9184 50568 0 _0625_
rlabel metal2 14280 50960 14280 50960 0 _0626_
rlabel metal2 7448 49672 7448 49672 0 _0627_
rlabel metal2 8232 50904 8232 50904 0 _0628_
rlabel metal2 10696 52976 10696 52976 0 _0629_
rlabel metal2 26488 55440 26488 55440 0 _0630_
rlabel metal2 29568 51912 29568 51912 0 _0631_
rlabel metal3 7000 39592 7000 39592 0 _0632_
rlabel metal2 7896 38920 7896 38920 0 _0633_
rlabel metal2 12376 43792 12376 43792 0 _0634_
rlabel metal2 15624 37072 15624 37072 0 _0635_
rlabel metal3 20048 42840 20048 42840 0 _0636_
rlabel metal2 24696 46592 24696 46592 0 _0637_
rlabel metal2 29624 52920 29624 52920 0 _0638_
rlabel metal2 24136 47320 24136 47320 0 _0639_
rlabel metal2 15512 36232 15512 36232 0 _0640_
rlabel metal2 19320 39984 19320 39984 0 _0641_
rlabel metal2 17416 41272 17416 41272 0 _0642_
rlabel metal2 11928 39312 11928 39312 0 _0643_
rlabel metal2 15848 39984 15848 39984 0 _0644_
rlabel metal2 22120 43792 22120 43792 0 _0645_
rlabel metal3 31416 47320 31416 47320 0 _0646_
rlabel metal2 16856 50120 16856 50120 0 _0647_
rlabel metal2 16968 39536 16968 39536 0 _0648_
rlabel metal2 24136 38920 24136 38920 0 _0649_
rlabel metal2 23352 48720 23352 48720 0 _0650_
rlabel metal2 15400 36064 15400 36064 0 _0651_
rlabel metal2 24248 35504 24248 35504 0 _0652_
rlabel metal3 25592 34888 25592 34888 0 _0653_
rlabel metal2 31640 50064 31640 50064 0 _0654_
rlabel metal2 26712 55328 26712 55328 0 _0655_
rlabel metal3 33208 50344 33208 50344 0 _0656_
rlabel metal2 34104 54208 34104 54208 0 _0657_
rlabel metal2 12488 53088 12488 53088 0 _0658_
rlabel metal2 26824 48048 26824 48048 0 _0659_
rlabel metal2 26544 49896 26544 49896 0 _0660_
rlabel metal2 10808 40208 10808 40208 0 _0661_
rlabel metal2 11480 38808 11480 38808 0 _0662_
rlabel metal2 26488 44240 26488 44240 0 _0663_
rlabel metal2 23800 39648 23800 39648 0 _0664_
rlabel metal3 24808 44296 24808 44296 0 _0665_
rlabel metal2 26320 47544 26320 47544 0 _0666_
rlabel metal2 33656 54656 33656 54656 0 _0667_
rlabel metal2 41832 54880 41832 54880 0 _0668_
rlabel metal2 48496 50456 48496 50456 0 _0669_
rlabel metal2 46200 51912 46200 51912 0 _0670_
rlabel metal2 48440 46984 48440 46984 0 _0671_
rlabel metal2 41496 53144 41496 53144 0 _0672_
rlabel metal2 18144 35000 18144 35000 0 _0673_
rlabel metal2 22456 54936 22456 54936 0 _0674_
rlabel metal2 12152 36344 12152 36344 0 _0675_
rlabel metal2 13608 50736 13608 50736 0 _0676_
rlabel metal2 8008 41328 8008 41328 0 _0677_
rlabel metal2 7336 41888 7336 41888 0 _0678_
rlabel metal2 11480 42728 11480 42728 0 _0679_
rlabel metal3 14140 53928 14140 53928 0 _0680_
rlabel metal3 13160 41944 13160 41944 0 _0681_
rlabel metal2 17192 36176 17192 36176 0 _0682_
rlabel metal2 12936 54208 12936 54208 0 _0683_
rlabel metal2 6552 52276 6552 52276 0 _0684_
rlabel metal2 19656 53872 19656 53872 0 _0685_
rlabel metal3 20328 53928 20328 53928 0 _0686_
rlabel metal2 8120 45696 8120 45696 0 _0687_
rlabel metal2 18144 43512 18144 43512 0 _0688_
rlabel metal2 18200 44968 18200 44968 0 _0689_
rlabel metal2 20496 45752 20496 45752 0 _0690_
rlabel metal2 11256 46032 11256 46032 0 _0691_
rlabel metal2 9240 39312 9240 39312 0 _0692_
rlabel metal2 19768 41664 19768 41664 0 _0693_
rlabel metal2 18760 46032 18760 46032 0 _0694_
rlabel metal2 19096 55776 19096 55776 0 _0695_
rlabel metal2 18424 54768 18424 54768 0 _0696_
rlabel metal2 12376 52360 12376 52360 0 _0697_
rlabel metal2 12824 54712 12824 54712 0 _0698_
rlabel metal2 17528 54768 17528 54768 0 _0699_
rlabel metal2 39032 53200 39032 53200 0 _0700_
rlabel metal3 48384 47992 48384 47992 0 _0701_
rlabel metal2 47152 51576 47152 51576 0 _0702_
rlabel metal2 24360 46088 24360 46088 0 _0703_
rlabel metal2 20664 51128 20664 51128 0 _0704_
rlabel metal3 39872 53144 39872 53144 0 _0705_
rlabel metal2 25872 50232 25872 50232 0 _0706_
rlabel metal3 17528 41048 17528 41048 0 _0707_
rlabel metal2 17864 39200 17864 39200 0 _0708_
rlabel metal2 14168 52080 14168 52080 0 _0709_
rlabel metal2 21672 40600 21672 40600 0 _0710_
rlabel metal3 14392 35896 14392 35896 0 _0711_
rlabel metal2 22456 40320 22456 40320 0 _0712_
rlabel metal3 18088 35896 18088 35896 0 _0713_
rlabel metal2 26544 41048 26544 41048 0 _0714_
rlabel metal4 22232 41384 22232 41384 0 _0715_
rlabel metal3 10808 40376 10808 40376 0 _0716_
rlabel metal2 10584 41048 10584 41048 0 _0717_
rlabel metal2 15288 43624 15288 43624 0 _0718_
rlabel metal2 17752 43624 17752 43624 0 _0719_
rlabel metal2 12432 50680 12432 50680 0 _0720_
rlabel metal4 20776 51912 20776 51912 0 _0721_
rlabel metal2 20440 51688 20440 51688 0 _0722_
rlabel metal3 23128 52136 23128 52136 0 _0723_
rlabel metal3 39200 53032 39200 53032 0 _0724_
rlabel metal3 41384 53928 41384 53928 0 _0725_
rlabel metal3 40432 53816 40432 53816 0 _0726_
rlabel metal3 40880 53592 40880 53592 0 _0727_
rlabel metal2 41272 54544 41272 54544 0 _0728_
rlabel metal2 41216 55160 41216 55160 0 _0729_
rlabel metal2 48048 45976 48048 45976 0 _0730_
rlabel metal2 49280 54376 49280 54376 0 _0731_
rlabel metal2 30632 49560 30632 49560 0 _0732_
rlabel metal2 35784 49252 35784 49252 0 _0733_
rlabel metal2 25928 45304 25928 45304 0 _0734_
rlabel metal3 19488 42056 19488 42056 0 _0735_
rlabel metal2 19880 47600 19880 47600 0 _0736_
rlabel metal2 27720 54768 27720 54768 0 _0737_
rlabel metal3 29512 53480 29512 53480 0 _0738_
rlabel metal2 23240 43512 23240 43512 0 _0739_
rlabel metal2 17976 47264 17976 47264 0 _0740_
rlabel metal4 27272 49112 27272 49112 0 _0741_
rlabel metal2 12432 54376 12432 54376 0 _0742_
rlabel metal2 27832 50512 27832 50512 0 _0743_
rlabel metal2 29792 51688 29792 51688 0 _0744_
rlabel metal3 19208 55776 19208 55776 0 _0745_
rlabel metal3 18256 42616 18256 42616 0 _0746_
rlabel metal3 21056 49672 21056 49672 0 _0747_
rlabel metal2 18760 49952 18760 49952 0 _0748_
rlabel metal3 25760 54488 25760 54488 0 _0749_
rlabel metal3 40992 54488 40992 54488 0 _0750_
rlabel metal2 44968 54320 44968 54320 0 _0751_
rlabel metal2 38976 55048 38976 55048 0 _0752_
rlabel metal2 36008 55328 36008 55328 0 _0753_
rlabel metal2 24136 49168 24136 49168 0 _0754_
rlabel metal2 23240 47208 23240 47208 0 _0755_
rlabel metal3 20944 50568 20944 50568 0 _0756_
rlabel metal3 23072 51128 23072 51128 0 _0757_
rlabel metal3 23408 49896 23408 49896 0 _0758_
rlabel metal2 9800 45472 9800 45472 0 _0759_
rlabel metal2 19992 45136 19992 45136 0 _0760_
rlabel metal2 20328 43512 20328 43512 0 _0761_
rlabel metal2 14728 43904 14728 43904 0 _0762_
rlabel metal2 23576 45528 23576 45528 0 _0763_
rlabel metal2 15176 41216 15176 41216 0 _0764_
rlabel metal3 16912 43400 16912 43400 0 _0765_
rlabel metal2 18424 43568 18424 43568 0 _0766_
rlabel metal3 24640 50344 24640 50344 0 _0767_
rlabel metal2 26824 49336 26824 49336 0 _0768_
rlabel metal3 42952 55272 42952 55272 0 _0769_
rlabel metal3 20944 48216 20944 48216 0 _0770_
rlabel metal2 21112 56784 21112 56784 0 _0771_
rlabel metal2 22400 41160 22400 41160 0 _0772_
rlabel metal2 24304 53480 24304 53480 0 _0773_
rlabel metal2 18760 33824 18760 33824 0 _0774_
rlabel metal2 19096 34328 19096 34328 0 _0775_
rlabel metal2 28504 54040 28504 54040 0 _0776_
rlabel metal2 13384 53984 13384 53984 0 _0777_
rlabel metal2 12264 50904 12264 50904 0 _0778_
rlabel metal2 14112 50792 14112 50792 0 _0779_
rlabel metal2 15736 51128 15736 51128 0 _0780_
rlabel metal2 25368 39928 25368 39928 0 _0781_
rlabel metal2 14392 52192 14392 52192 0 _0782_
rlabel metal3 18424 52248 18424 52248 0 _0783_
rlabel metal2 22792 54376 22792 54376 0 _0784_
rlabel metal2 28392 54768 28392 54768 0 _0785_
rlabel metal3 39256 54376 39256 54376 0 _0786_
rlabel metal3 40656 53704 40656 53704 0 _0787_
rlabel metal2 45640 51520 45640 51520 0 _0788_
rlabel metal2 44296 48832 44296 48832 0 _0789_
rlabel metal3 12208 38920 12208 38920 0 _0790_
rlabel metal2 16296 43400 16296 43400 0 _0791_
rlabel metal2 16632 45080 16632 45080 0 _0792_
rlabel metal2 21336 46984 21336 46984 0 _0793_
rlabel metal3 19208 50344 19208 50344 0 _0794_
rlabel metal2 18312 47376 18312 47376 0 _0795_
rlabel metal3 20104 51072 20104 51072 0 _0796_
rlabel metal2 18144 46872 18144 46872 0 _0797_
rlabel metal2 21224 34440 21224 34440 0 _0798_
rlabel metal2 31752 51072 31752 51072 0 _0799_
rlabel metal3 31584 53704 31584 53704 0 _0800_
rlabel metal3 31024 46984 31024 46984 0 _0801_
rlabel metal2 39480 52192 39480 52192 0 _0802_
rlabel metal3 40712 52136 40712 52136 0 _0803_
rlabel metal2 43456 51240 43456 51240 0 _0804_
rlabel metal2 37576 51352 37576 51352 0 _0805_
rlabel metal2 21392 41048 21392 41048 0 _0806_
rlabel metal3 24192 42728 24192 42728 0 _0807_
rlabel metal2 32088 39368 32088 39368 0 _0808_
rlabel metal2 24024 36400 24024 36400 0 _0809_
rlabel metal2 15400 40432 15400 40432 0 _0810_
rlabel metal2 18088 47264 18088 47264 0 _0811_
rlabel metal3 23688 38696 23688 38696 0 _0812_
rlabel metal2 22120 36792 22120 36792 0 _0813_
rlabel metal2 22792 36400 22792 36400 0 _0814_
rlabel metal2 24360 36120 24360 36120 0 _0815_
rlabel metal3 17248 48664 17248 48664 0 _0816_
rlabel metal2 25648 48888 25648 48888 0 _0817_
rlabel metal3 19824 48440 19824 48440 0 _0818_
rlabel metal2 27944 45528 27944 45528 0 _0819_
rlabel metal2 21896 37856 21896 37856 0 _0820_
rlabel metal2 34552 44688 34552 44688 0 _0821_
rlabel metal2 35336 47488 35336 47488 0 _0822_
rlabel metal2 34664 44184 34664 44184 0 _0823_
rlabel metal2 31472 51576 31472 51576 0 _0824_
rlabel metal2 22344 51688 22344 51688 0 _0825_
rlabel metal2 19096 44912 19096 44912 0 _0826_
rlabel metal2 30968 51016 30968 51016 0 _0827_
rlabel metal2 38808 50428 38808 50428 0 _0828_
rlabel metal3 30464 50792 30464 50792 0 _0829_
rlabel metal3 34664 50792 34664 50792 0 _0830_
rlabel metal2 41272 52248 41272 52248 0 _0831_
rlabel metal2 42504 53032 42504 53032 0 _0832_
rlabel metal2 42840 54208 42840 54208 0 _0833_
rlabel metal2 43400 54600 43400 54600 0 _0834_
rlabel metal2 43848 54824 43848 54824 0 _0835_
rlabel metal2 44520 55272 44520 55272 0 _0836_
rlabel metal2 50792 54656 50792 54656 0 _0837_
rlabel metal2 48216 55104 48216 55104 0 _0838_
rlabel metal2 35560 54040 35560 54040 0 _0839_
rlabel metal2 37240 54432 37240 54432 0 _0840_
rlabel metal2 36680 54768 36680 54768 0 _0841_
rlabel metal3 28056 47264 28056 47264 0 _0842_
rlabel metal2 29344 49000 29344 49000 0 _0843_
rlabel metal2 23240 48104 23240 48104 0 _0844_
rlabel metal2 25592 50848 25592 50848 0 _0845_
rlabel metal2 33768 51464 33768 51464 0 _0846_
rlabel metal2 24024 39200 24024 39200 0 _0847_
rlabel metal2 12376 47992 12376 47992 0 _0848_
rlabel metal2 23800 44856 23800 44856 0 _0849_
rlabel metal2 24808 46032 24808 46032 0 _0850_
rlabel metal2 13776 50792 13776 50792 0 _0851_
rlabel metal2 15960 47992 15960 47992 0 _0852_
rlabel metal3 22344 45192 22344 45192 0 _0853_
rlabel via2 23016 44296 23016 44296 0 _0854_
rlabel metal2 17752 44744 17752 44744 0 _0855_
rlabel metal2 24024 44744 24024 44744 0 _0856_
rlabel metal3 25144 45192 25144 45192 0 _0857_
rlabel metal2 25816 46312 25816 46312 0 _0858_
rlabel metal2 34888 52024 34888 52024 0 _0859_
rlabel metal2 36120 53424 36120 53424 0 _0860_
rlabel metal2 46424 54544 46424 54544 0 _0861_
rlabel metal3 49224 52248 49224 52248 0 _0862_
rlabel metal2 41664 47320 41664 47320 0 _0863_
rlabel metal2 40936 48664 40936 48664 0 _0864_
rlabel metal2 41048 48720 41048 48720 0 _0865_
rlabel metal2 10920 48664 10920 48664 0 _0866_
rlabel metal3 16184 43400 16184 43400 0 _0867_
rlabel metal2 13496 47712 13496 47712 0 _0868_
rlabel metal2 14952 43568 14952 43568 0 _0869_
rlabel metal2 13944 46424 13944 46424 0 _0870_
rlabel metal3 12600 49000 12600 49000 0 _0871_
rlabel metal2 14056 48104 14056 48104 0 _0872_
rlabel metal2 15064 53144 15064 53144 0 _0873_
rlabel metal2 20608 34216 20608 34216 0 _0874_
rlabel metal2 37016 40824 37016 40824 0 _0875_
rlabel metal2 19152 40600 19152 40600 0 _0876_
rlabel metal2 37912 46760 37912 46760 0 _0877_
rlabel metal2 39928 48552 39928 48552 0 _0878_
rlabel metal2 39368 34160 39368 34160 0 _0879_
rlabel metal3 40656 43512 40656 43512 0 _0880_
rlabel metal2 40152 48720 40152 48720 0 _0881_
rlabel metal2 45864 51576 45864 51576 0 _0882_
rlabel metal2 42728 51688 42728 51688 0 _0883_
rlabel metal2 43792 51128 43792 51128 0 _0884_
rlabel metal2 44072 51632 44072 51632 0 _0885_
rlabel metal2 20328 50736 20328 50736 0 _0886_
rlabel metal2 21672 50064 21672 50064 0 _0887_
rlabel metal2 28392 51072 28392 51072 0 _0888_
rlabel metal2 24696 35952 24696 35952 0 _0889_
rlabel metal2 21672 41160 21672 41160 0 _0890_
rlabel metal2 22792 42224 22792 42224 0 _0891_
rlabel metal2 22456 46256 22456 46256 0 _0892_
rlabel metal3 21672 39816 21672 39816 0 _0893_
rlabel metal2 21896 46592 21896 46592 0 _0894_
rlabel metal2 16744 44800 16744 44800 0 _0895_
rlabel metal3 21000 46648 21000 46648 0 _0896_
rlabel metal2 24024 46592 24024 46592 0 _0897_
rlabel metal2 42504 51128 42504 51128 0 _0898_
rlabel metal3 44632 52248 44632 52248 0 _0899_
rlabel metal3 44240 52136 44240 52136 0 _0900_
rlabel metal2 45752 52472 45752 52472 0 _0901_
rlabel metal2 47768 53760 47768 53760 0 _0902_
rlabel metal2 50008 54936 50008 54936 0 _0903_
rlabel metal2 51464 54488 51464 54488 0 _0904_
rlabel metal2 52416 55160 52416 55160 0 _0905_
rlabel metal2 45864 53032 45864 53032 0 _0906_
rlabel metal2 50120 53256 50120 53256 0 _0907_
rlabel metal2 37240 52808 37240 52808 0 _0908_
rlabel metal3 36064 49784 36064 49784 0 _0909_
rlabel metal2 16184 45472 16184 45472 0 _0910_
rlabel metal2 18536 49280 18536 49280 0 _0911_
rlabel metal2 29176 49056 29176 49056 0 _0912_
rlabel metal2 25592 47880 25592 47880 0 _0913_
rlabel metal2 27720 45640 27720 45640 0 _0914_
rlabel metal2 27608 48552 27608 48552 0 _0915_
rlabel metal2 27720 48272 27720 48272 0 _0916_
rlabel metal2 28056 48216 28056 48216 0 _0917_
rlabel metal2 29512 49392 29512 49392 0 _0918_
rlabel metal3 26740 40600 26740 40600 0 _0919_
rlabel metal3 32032 48776 32032 48776 0 _0920_
rlabel metal2 32760 49112 32760 49112 0 _0921_
rlabel metal2 33880 49672 33880 49672 0 _0922_
rlabel metal2 38472 51072 38472 51072 0 _0923_
rlabel metal2 48664 51408 48664 51408 0 _0924_
rlabel metal2 46368 49896 46368 49896 0 _0925_
rlabel metal2 11032 49448 11032 49448 0 _0926_
rlabel metal2 10360 44016 10360 44016 0 _0927_
rlabel metal4 12040 43624 12040 43624 0 _0928_
rlabel metal2 11704 47264 11704 47264 0 _0929_
rlabel metal2 19208 49168 19208 49168 0 _0930_
rlabel metal2 16296 49336 16296 49336 0 _0931_
rlabel metal3 22232 34888 22232 34888 0 _0932_
rlabel metal4 25256 39760 25256 39760 0 _0933_
rlabel metal2 14616 47880 14616 47880 0 _0934_
rlabel metal2 17528 45752 17528 45752 0 _0935_
rlabel metal2 18424 41440 18424 41440 0 _0936_
rlabel metal2 16968 46704 16968 46704 0 _0937_
rlabel metal2 16856 49056 16856 49056 0 _0938_
rlabel metal3 46704 49000 46704 49000 0 _0939_
rlabel metal2 43736 49896 43736 49896 0 _0940_
rlabel metal3 45136 50456 45136 50456 0 _0941_
rlabel metal2 40488 42952 40488 42952 0 _0942_
rlabel metal2 22344 46424 22344 46424 0 _0943_
rlabel metal2 22456 48328 22456 48328 0 _0944_
rlabel metal2 23016 49448 23016 49448 0 _0945_
rlabel metal2 18648 47880 18648 47880 0 _0946_
rlabel metal3 17696 46872 17696 46872 0 _0947_
rlabel metal3 20720 45752 20720 45752 0 _0948_
rlabel metal2 19264 47656 19264 47656 0 _0949_
rlabel metal3 37352 47432 37352 47432 0 _0950_
rlabel metal2 39032 49504 39032 49504 0 _0951_
rlabel metal2 39816 49392 39816 49392 0 _0952_
rlabel metal3 43568 49784 43568 49784 0 _0953_
rlabel metal2 48888 50512 48888 50512 0 _0954_
rlabel metal3 48216 50568 48216 50568 0 _0955_
rlabel metal2 50680 50624 50680 50624 0 _0956_
rlabel metal3 49952 52136 49952 52136 0 _0957_
rlabel metal2 51352 53144 51352 53144 0 _0958_
rlabel metal3 48664 54488 48664 54488 0 _0959_
rlabel metal2 46872 54208 46872 54208 0 _0960_
rlabel metal3 48048 54600 48048 54600 0 _0961_
rlabel metal3 52640 54488 52640 54488 0 _0962_
rlabel metal2 52808 53312 52808 53312 0 _0963_
rlabel metal2 53480 53312 53480 53312 0 _0964_
rlabel metal3 50512 50456 50512 50456 0 _0965_
rlabel metal2 51016 49616 51016 49616 0 _0966_
rlabel metal3 29064 45192 29064 45192 0 _0967_
rlabel metal2 29792 35672 29792 35672 0 _0968_
rlabel metal2 26264 37800 26264 37800 0 _0969_
rlabel metal2 28224 40600 28224 40600 0 _0970_
rlabel metal3 24136 40936 24136 40936 0 _0971_
rlabel metal3 26292 41832 26292 41832 0 _0972_
rlabel metal2 27944 42280 27944 42280 0 _0973_
rlabel metal2 33656 41440 33656 41440 0 _0974_
rlabel metal2 27720 40376 27720 40376 0 _0975_
rlabel metal2 30072 45080 30072 45080 0 _0976_
rlabel metal2 29848 42952 29848 42952 0 _0977_
rlabel metal2 29288 42224 29288 42224 0 _0978_
rlabel metal2 30184 42616 30184 42616 0 _0979_
rlabel metal3 33600 43512 33600 43512 0 _0980_
rlabel metal2 37352 51408 37352 51408 0 _0981_
rlabel metal2 36624 43624 36624 43624 0 _0982_
rlabel metal2 38472 43120 38472 43120 0 _0983_
rlabel metal2 50232 45192 50232 45192 0 _0984_
rlabel metal2 45136 46648 45136 46648 0 _0985_
rlabel metal2 45528 48496 45528 48496 0 _0986_
rlabel metal2 21448 50120 21448 50120 0 _0987_
rlabel metal2 17640 45696 17640 45696 0 _0988_
rlabel metal2 19096 42560 19096 42560 0 _0989_
rlabel metal2 13384 45304 13384 45304 0 _0990_
rlabel metal2 15736 45976 15736 45976 0 _0991_
rlabel metal2 16408 46592 16408 46592 0 _0992_
rlabel metal2 22848 50008 22848 50008 0 _0993_
rlabel metal3 45528 48216 45528 48216 0 _0994_
rlabel metal3 46592 47432 46592 47432 0 _0995_
rlabel metal2 50792 47488 50792 47488 0 _0996_
rlabel metal2 40824 47712 40824 47712 0 _0997_
rlabel metal2 42280 41272 42280 41272 0 _0998_
rlabel metal2 23016 42392 23016 42392 0 _0999_
rlabel metal3 22008 43400 22008 43400 0 _1000_
rlabel metal2 24136 42448 24136 42448 0 _1001_
rlabel metal3 22120 41664 22120 41664 0 _1002_
rlabel metal2 22344 41552 22344 41552 0 _1003_
rlabel metal2 21672 42336 21672 42336 0 _1004_
rlabel metal2 21448 41664 21448 41664 0 _1005_
rlabel metal2 21560 42224 21560 42224 0 _1006_
rlabel metal2 39368 43848 39368 43848 0 _1007_
rlabel metal2 39256 44912 39256 44912 0 _1008_
rlabel metal2 48776 46928 48776 46928 0 _1009_
rlabel metal2 49112 47488 49112 47488 0 _1010_
rlabel metal2 50456 47432 50456 47432 0 _1011_
rlabel metal2 49840 47992 49840 47992 0 _1012_
rlabel metal2 50904 49000 50904 49000 0 _1013_
rlabel metal2 53928 50176 53928 50176 0 _1014_
rlabel via2 52360 50680 52360 50680 0 _1015_
rlabel metal2 50904 53760 50904 53760 0 _1016_
rlabel metal2 52920 52584 52920 52584 0 _1017_
rlabel metal2 53480 50680 53480 50680 0 _1018_
rlabel metal2 54600 51016 54600 51016 0 _1019_
rlabel metal2 52248 46928 52248 46928 0 _1020_
rlabel metal2 52024 46872 52024 46872 0 _1021_
rlabel metal2 53144 47768 53144 47768 0 _1022_
rlabel metal2 31528 42280 31528 42280 0 _1023_
rlabel metal2 27384 45696 27384 45696 0 _1024_
rlabel metal2 31080 43960 31080 43960 0 _1025_
rlabel metal3 30184 44296 30184 44296 0 _1026_
rlabel metal2 26600 43176 26600 43176 0 _1027_
rlabel metal2 30968 44184 30968 44184 0 _1028_
rlabel metal2 34328 39480 34328 39480 0 _1029_
rlabel metal2 36792 43904 36792 43904 0 _1030_
rlabel metal2 37632 39592 37632 39592 0 _1031_
rlabel metal2 37856 42840 37856 42840 0 _1032_
rlabel metal2 50680 44352 50680 44352 0 _1033_
rlabel metal2 45528 46872 45528 46872 0 _1034_
rlabel metal2 20328 46368 20328 46368 0 _1035_
rlabel metal2 20384 45976 20384 45976 0 _1036_
rlabel metal2 21560 45528 21560 45528 0 _1037_
rlabel metal2 20104 35168 20104 35168 0 _1038_
rlabel metal3 36176 42280 36176 42280 0 _1039_
rlabel metal2 36008 44688 36008 44688 0 _1040_
rlabel metal2 43512 44688 43512 44688 0 _1041_
rlabel metal2 46872 45136 46872 45136 0 _1042_
rlabel metal3 46256 45080 46256 45080 0 _1043_
rlabel metal2 41272 44632 41272 44632 0 _1044_
rlabel metal2 38584 46536 38584 46536 0 _1045_
rlabel metal3 30856 47656 30856 47656 0 _1046_
rlabel metal3 30520 47544 30520 47544 0 _1047_
rlabel metal3 33768 47656 33768 47656 0 _1048_
rlabel metal2 19320 44632 19320 44632 0 _1049_
rlabel metal3 31528 47432 31528 47432 0 _1050_
rlabel metal3 25788 47544 25788 47544 0 _1051_
rlabel metal2 35000 47488 35000 47488 0 _1052_
rlabel metal2 35728 46760 35728 46760 0 _1053_
rlabel metal2 35560 47544 35560 47544 0 _1054_
rlabel metal3 39648 45752 39648 45752 0 _1055_
rlabel metal2 39816 43792 39816 43792 0 _1056_
rlabel metal2 42504 41608 42504 41608 0 _1057_
rlabel metal2 35112 47096 35112 47096 0 _1058_
rlabel metal2 39928 46704 39928 46704 0 _1059_
rlabel metal2 41048 44520 41048 44520 0 _1060_
rlabel metal2 40824 44576 40824 44576 0 _1061_
rlabel metal3 44464 44520 44464 44520 0 _1062_
rlabel metal3 48384 45192 48384 45192 0 _1063_
rlabel metal2 47432 44800 47432 44800 0 _1064_
rlabel metal2 50848 44408 50848 44408 0 _1065_
rlabel metal2 51800 45528 51800 45528 0 _1066_
rlabel metal2 54264 49448 54264 49448 0 _1067_
rlabel metal2 52808 47768 52808 47768 0 _1068_
rlabel metal3 53536 49112 53536 49112 0 _1069_
rlabel metal2 54712 49728 54712 49728 0 _1070_
rlabel metal2 52248 43568 52248 43568 0 _1071_
rlabel metal2 37800 39816 37800 39816 0 _1072_
rlabel metal2 38808 36232 38808 36232 0 _1073_
rlabel metal2 31192 40320 31192 40320 0 _1074_
rlabel metal2 23688 39116 23688 39116 0 _1075_
rlabel metal2 25032 39928 25032 39928 0 _1076_
rlabel metal2 31192 42000 31192 42000 0 _1077_
rlabel metal3 28504 38808 28504 38808 0 _1078_
rlabel metal2 35112 41216 35112 41216 0 _1079_
rlabel metal2 34664 41608 34664 41608 0 _1080_
rlabel metal3 36512 41832 36512 41832 0 _1081_
rlabel metal2 47880 41104 47880 41104 0 _1082_
rlabel metal2 45360 41944 45360 41944 0 _1083_
rlabel metal2 29680 38808 29680 38808 0 _1084_
rlabel metal2 29008 38024 29008 38024 0 _1085_
rlabel metal2 28056 41664 28056 41664 0 _1086_
rlabel metal2 28728 39620 28728 39620 0 _1087_
rlabel metal2 28280 37688 28280 37688 0 _1088_
rlabel metal3 28952 38024 28952 38024 0 _1089_
rlabel metal2 29512 34888 29512 34888 0 _1090_
rlabel metal2 29288 36736 29288 36736 0 _1091_
rlabel metal2 44744 40264 44744 40264 0 _1092_
rlabel metal2 46424 41496 46424 41496 0 _1093_
rlabel metal2 41944 41216 41944 41216 0 _1094_
rlabel metal2 34440 44520 34440 44520 0 _1095_
rlabel metal2 34888 40880 34888 40880 0 _1096_
rlabel metal2 22400 39032 22400 39032 0 _1097_
rlabel metal3 22792 39704 22792 39704 0 _1098_
rlabel metal3 24248 38808 24248 38808 0 _1099_
rlabel metal3 23800 39592 23800 39592 0 _1100_
rlabel metal2 35896 40040 35896 40040 0 _1101_
rlabel metal2 38808 40768 38808 40768 0 _1102_
rlabel metal3 40712 41160 40712 41160 0 _1103_
rlabel metal3 43120 42616 43120 42616 0 _1104_
rlabel metal2 42168 41272 42168 41272 0 _1105_
rlabel metal2 45640 40880 45640 40880 0 _1106_
rlabel metal3 47376 41272 47376 41272 0 _1107_
rlabel metal3 46536 41944 46536 41944 0 _1108_
rlabel metal2 41160 41160 41160 41160 0 _1109_
rlabel metal3 44576 41384 44576 41384 0 _1110_
rlabel metal2 48440 42392 48440 42392 0 _1111_
rlabel metal2 51576 42336 51576 42336 0 _1112_
rlabel metal2 51352 42728 51352 42728 0 _1113_
rlabel metal2 52360 43456 52360 43456 0 _1114_
rlabel metal2 54544 45080 54544 45080 0 _1115_
rlabel metal2 53928 45304 53928 45304 0 _1116_
rlabel metal2 52584 47376 52584 47376 0 _1117_
rlabel metal3 52976 46648 52976 46648 0 _1118_
rlabel metal2 53648 45192 53648 45192 0 _1119_
rlabel metal2 54152 44968 54152 44968 0 _1120_
rlabel metal2 55440 45080 55440 45080 0 _1121_
rlabel metal2 47096 36512 47096 36512 0 _1122_
rlabel metal2 47320 41552 47320 41552 0 _1123_
rlabel metal2 51016 40768 51016 40768 0 _1124_
rlabel metal3 35336 38920 35336 38920 0 _1125_
rlabel metal2 32088 36792 32088 36792 0 _1126_
rlabel metal2 29680 35896 29680 35896 0 _1127_
rlabel metal2 34888 37688 34888 37688 0 _1128_
rlabel metal3 34664 39592 34664 39592 0 _1129_
rlabel metal3 35056 37800 35056 37800 0 _1130_
rlabel metal2 35840 35672 35840 35672 0 _1131_
rlabel metal3 37016 38696 37016 38696 0 _1132_
rlabel metal3 44016 38696 44016 38696 0 _1133_
rlabel metal2 30072 37464 30072 37464 0 _1134_
rlabel metal2 31528 38920 31528 38920 0 _1135_
rlabel metal3 26740 36568 26740 36568 0 _1136_
rlabel metal2 26712 37520 26712 37520 0 _1137_
rlabel metal2 31808 40488 31808 40488 0 _1138_
rlabel metal2 32088 39816 32088 39816 0 _1139_
rlabel metal3 27608 40936 27608 40936 0 _1140_
rlabel metal3 42728 38808 42728 38808 0 _1141_
rlabel metal2 45976 39144 45976 39144 0 _1142_
rlabel metal3 44128 38920 44128 38920 0 _1143_
rlabel metal2 44800 39368 44800 39368 0 _1144_
rlabel metal3 28952 39368 28952 39368 0 _1145_
rlabel metal2 28504 40320 28504 40320 0 _1146_
rlabel metal3 44576 37464 44576 37464 0 _1147_
rlabel metal3 45808 38808 45808 38808 0 _1148_
rlabel metal2 46312 39144 46312 39144 0 _1149_
rlabel metal2 49000 38920 49000 38920 0 _1150_
rlabel metal2 48664 39480 48664 39480 0 _1151_
rlabel metal3 47264 39592 47264 39592 0 _1152_
rlabel metal3 49336 39816 49336 39816 0 _1153_
rlabel metal2 51128 39312 51128 39312 0 _1154_
rlabel metal2 51800 40488 51800 40488 0 _1155_
rlabel metal2 52136 40880 52136 40880 0 _1156_
rlabel metal3 52416 41048 52416 41048 0 _1157_
rlabel metal2 54936 43932 54936 43932 0 _1158_
rlabel metal3 53032 42168 53032 42168 0 _1159_
rlabel metal2 54320 43400 54320 43400 0 _1160_
rlabel metal3 56168 43512 56168 43512 0 _1161_
rlabel metal2 53480 40768 53480 40768 0 _1162_
rlabel metal2 51296 40152 51296 40152 0 _1163_
rlabel metal2 53368 40600 53368 40600 0 _1164_
rlabel metal2 54488 40768 54488 40768 0 _1165_
rlabel metal3 53872 44296 53872 44296 0 _1166_
rlabel metal2 54656 41160 54656 41160 0 _1167_
rlabel metal2 53256 39256 53256 39256 0 _1168_
rlabel metal2 29512 46368 29512 46368 0 _1169_
rlabel metal2 30632 45472 30632 45472 0 _1170_
rlabel metal2 29624 44856 29624 44856 0 _1171_
rlabel metal3 30016 45080 30016 45080 0 _1172_
rlabel metal2 31304 45584 31304 45584 0 _1173_
rlabel metal2 42168 45584 42168 45584 0 _1174_
rlabel metal2 41384 45360 41384 45360 0 _1175_
rlabel metal3 42224 43512 42224 43512 0 _1176_
rlabel metal2 42952 43176 42952 43176 0 _1177_
rlabel metal3 47376 42728 47376 42728 0 _1178_
rlabel metal2 44912 44296 44912 44296 0 _1179_
rlabel metal3 32144 42728 32144 42728 0 _1180_
rlabel metal3 34160 42616 34160 42616 0 _1181_
rlabel metal3 34832 39704 34832 39704 0 _1182_
rlabel metal2 45416 42896 45416 42896 0 _1183_
rlabel metal3 44184 44072 44184 44072 0 _1184_
rlabel metal2 44968 43400 44968 43400 0 _1185_
rlabel metal2 49448 43120 49448 43120 0 _1186_
rlabel metal2 49336 42952 49336 42952 0 _1187_
rlabel metal2 51072 38024 51072 38024 0 _1188_
rlabel metal3 36792 37352 36792 37352 0 _1189_
rlabel metal2 27944 36568 27944 36568 0 _1190_
rlabel metal2 25368 37576 25368 37576 0 _1191_
rlabel metal3 33040 37912 33040 37912 0 _1192_
rlabel metal2 39032 37520 39032 37520 0 _1193_
rlabel metal3 44576 37352 44576 37352 0 _1194_
rlabel metal2 51464 37352 51464 37352 0 _1195_
rlabel metal3 52528 38808 52528 38808 0 _1196_
rlabel metal2 55160 39648 55160 39648 0 _1197_
rlabel metal2 55272 40488 55272 40488 0 _1198_
rlabel metal2 55048 40600 55048 40600 0 _1199_
rlabel metal2 50512 37464 50512 37464 0 _1200_
rlabel metal2 50960 37240 50960 37240 0 _1201_
rlabel metal2 26152 33320 26152 33320 0 _1202_
rlabel metal2 25592 35224 25592 35224 0 _1203_
rlabel metal2 32872 34384 32872 34384 0 _1204_
rlabel metal2 38696 35448 38696 35448 0 _1205_
rlabel metal2 38360 35952 38360 35952 0 _1206_
rlabel metal3 44296 35672 44296 35672 0 _1207_
rlabel metal2 32424 36736 32424 36736 0 _1208_
rlabel metal2 31416 36512 31416 36512 0 _1209_
rlabel metal3 34552 37576 34552 37576 0 _1210_
rlabel metal2 41048 37464 41048 37464 0 _1211_
rlabel metal2 41944 37240 41944 37240 0 _1212_
rlabel metal2 41384 37688 41384 37688 0 _1213_
rlabel metal2 47432 35784 47432 35784 0 _1214_
rlabel metal3 35056 36344 35056 36344 0 _1215_
rlabel metal2 44184 36960 44184 36960 0 _1216_
rlabel metal3 45136 37240 45136 37240 0 _1217_
rlabel metal2 47208 36176 47208 36176 0 _1218_
rlabel metal2 49560 36064 49560 36064 0 _1219_
rlabel metal3 51044 37352 51044 37352 0 _1220_
rlabel metal2 53928 37912 53928 37912 0 _1221_
rlabel metal2 53032 36400 53032 36400 0 _1222_
rlabel metal2 54264 38080 54264 38080 0 _1223_
rlabel metal2 54152 39760 54152 39760 0 _1224_
rlabel metal2 54376 37744 54376 37744 0 _1225_
rlabel metal2 55496 37632 55496 37632 0 _1226_
rlabel metal2 30408 35000 30408 35000 0 _1227_
rlabel metal2 32424 37912 32424 37912 0 _1228_
rlabel metal2 34328 33992 34328 33992 0 _1229_
rlabel metal2 47544 35000 47544 35000 0 _1230_
rlabel metal2 43624 32928 43624 32928 0 _1231_
rlabel metal3 45472 32648 45472 32648 0 _1232_
rlabel metal2 44856 35168 44856 35168 0 _1233_
rlabel metal2 44968 35728 44968 35728 0 _1234_
rlabel metal2 45976 35392 45976 35392 0 _1235_
rlabel metal3 47824 32760 47824 32760 0 _1236_
rlabel metal2 47992 32872 47992 32872 0 _1237_
rlabel metal2 48328 32200 48328 32200 0 _1238_
rlabel metal2 37240 35224 37240 35224 0 _1239_
rlabel metal3 36848 34888 36848 34888 0 _1240_
rlabel metal2 45192 34440 45192 34440 0 _1241_
rlabel metal2 48216 32592 48216 32592 0 _1242_
rlabel metal2 49784 32256 49784 32256 0 _1243_
rlabel metal3 49952 33208 49952 33208 0 _1244_
rlabel metal2 53032 34552 53032 34552 0 _1245_
rlabel metal2 47992 35224 47992 35224 0 _1246_
rlabel metal2 50568 34216 50568 34216 0 _1247_
rlabel metal3 53760 35672 53760 35672 0 _1248_
rlabel metal2 53816 36848 53816 36848 0 _1249_
rlabel metal2 53592 37296 53592 37296 0 _1250_
rlabel metal2 53424 35672 53424 35672 0 _1251_
rlabel metal2 54376 34944 54376 34944 0 _1252_
rlabel metal2 55216 34216 55216 34216 0 _1253_
rlabel metal2 30240 34888 30240 34888 0 _1254_
rlabel metal2 41272 36176 41272 36176 0 _1255_
rlabel metal2 41608 36176 41608 36176 0 _1256_
rlabel metal2 42728 35672 42728 35672 0 _1257_
rlabel metal3 6272 25368 6272 25368 0 _1258_
rlabel metal3 44912 34328 44912 34328 0 _1259_
rlabel metal3 47936 33320 47936 33320 0 _1260_
rlabel metal2 50904 33264 50904 33264 0 _1261_
rlabel metal2 50344 32984 50344 32984 0 _1262_
rlabel metal2 51912 33656 51912 33656 0 _1263_
rlabel metal2 52808 33936 52808 33936 0 _1264_
rlabel metal2 53872 33208 53872 33208 0 _1265_
rlabel metal2 46816 33880 46816 33880 0 _1266_
rlabel metal2 46424 34552 46424 34552 0 _1267_
rlabel metal2 5768 24416 5768 24416 0 _1268_
rlabel metal3 47824 34888 47824 34888 0 _1269_
rlabel metal2 52024 34552 52024 34552 0 _1270_
rlabel metal2 49224 34776 49224 34776 0 _1271_
rlabel metal3 50456 34104 50456 34104 0 _1272_
rlabel metal2 49336 33824 49336 33824 0 _1273_
rlabel metal2 49896 34552 49896 34552 0 _1274_
rlabel metal2 49616 34888 49616 34888 0 _1275_
rlabel metal2 46032 55160 46032 55160 0 _1276_
rlabel metal3 16352 18536 16352 18536 0 _1277_
rlabel metal2 28168 23576 28168 23576 0 _1278_
rlabel metal3 26712 14392 26712 14392 0 _1279_
rlabel metal2 28392 25088 28392 25088 0 _1280_
rlabel metal2 28168 22232 28168 22232 0 _1281_
rlabel metal2 9352 23520 9352 23520 0 _1282_
rlabel metal3 9296 20776 9296 20776 0 _1283_
rlabel metal2 11704 22792 11704 22792 0 _1284_
rlabel metal3 16520 10976 16520 10976 0 _1285_
rlabel metal2 8456 11536 8456 11536 0 _1286_
rlabel metal2 9800 18760 9800 18760 0 _1287_
rlabel metal3 14336 28616 14336 28616 0 _1288_
rlabel metal3 8680 11368 8680 11368 0 _1289_
rlabel metal3 9240 19208 9240 19208 0 _1290_
rlabel metal3 18648 26376 18648 26376 0 _1291_
rlabel metal2 15400 22624 15400 22624 0 _1292_
rlabel metal2 24024 19488 24024 19488 0 _1293_
rlabel metal3 11536 19880 11536 19880 0 _1294_
rlabel metal2 7896 18648 7896 18648 0 _1295_
rlabel metal2 19208 20160 19208 20160 0 _1296_
rlabel metal2 12992 20552 12992 20552 0 _1297_
rlabel metal2 11928 24248 11928 24248 0 _1298_
rlabel metal2 15064 18368 15064 18368 0 _1299_
rlabel via2 12936 24248 12936 24248 0 _1300_
rlabel metal2 13048 19432 13048 19432 0 _1301_
rlabel metal2 10640 25480 10640 25480 0 _1302_
rlabel metal2 11592 22064 11592 22064 0 _1303_
rlabel metal2 16632 20440 16632 20440 0 _1304_
rlabel metal3 7000 21560 7000 21560 0 _1305_
rlabel metal2 15400 19376 15400 19376 0 _1306_
rlabel metal2 12264 19992 12264 19992 0 _1307_
rlabel metal2 15848 20440 15848 20440 0 _1308_
rlabel metal2 17528 19600 17528 19600 0 _1309_
rlabel metal2 15848 18144 15848 18144 0 _1310_
rlabel metal2 18648 18200 18648 18200 0 _1311_
rlabel metal2 18088 22064 18088 22064 0 _1312_
rlabel metal2 18760 18816 18760 18816 0 _1313_
rlabel metal2 20160 18424 20160 18424 0 _1314_
rlabel metal2 21896 18928 21896 18928 0 _1315_
rlabel metal2 28504 18928 28504 18928 0 _1316_
rlabel metal3 26768 24584 26768 24584 0 _1317_
rlabel metal2 22792 14616 22792 14616 0 _1318_
rlabel metal3 26152 19320 26152 19320 0 _1319_
rlabel metal2 41608 21784 41608 21784 0 _1320_
rlabel metal2 5096 24752 5096 24752 0 _1321_
rlabel metal2 46200 24584 46200 24584 0 _1322_
rlabel metal2 40936 23520 40936 23520 0 _1323_
rlabel metal2 41496 23016 41496 23016 0 _1324_
rlabel metal2 17528 25424 17528 25424 0 _1325_
rlabel metal2 16184 25256 16184 25256 0 _1326_
rlabel metal2 15624 26208 15624 26208 0 _1327_
rlabel metal3 14448 26264 14448 26264 0 _1328_
rlabel metal3 16464 26264 16464 26264 0 _1329_
rlabel metal2 30968 24808 30968 24808 0 _1330_
rlabel metal3 19488 22344 19488 22344 0 _1331_
rlabel metal2 5096 17920 5096 17920 0 _1332_
rlabel metal2 29176 25536 29176 25536 0 _1333_
rlabel metal2 31192 24752 31192 24752 0 _1334_
rlabel metal2 8456 23520 8456 23520 0 _1335_
rlabel metal3 7336 19992 7336 19992 0 _1336_
rlabel metal2 9912 19264 9912 19264 0 _1337_
rlabel metal3 10024 23688 10024 23688 0 _1338_
rlabel metal2 20328 22792 20328 22792 0 _1339_
rlabel metal2 21448 19544 21448 19544 0 _1340_
rlabel metal2 22120 24024 22120 24024 0 _1341_
rlabel metal2 31528 23688 31528 23688 0 _1342_
rlabel metal2 8680 17808 8680 17808 0 _1343_
rlabel metal3 33544 24696 33544 24696 0 _1344_
rlabel metal2 42448 23912 42448 23912 0 _1345_
rlabel metal3 23576 25480 23576 25480 0 _1346_
rlabel metal2 23576 27664 23576 27664 0 _1347_
rlabel metal2 24472 23688 24472 23688 0 _1348_
rlabel metal2 17640 19936 17640 19936 0 _1349_
rlabel metal2 7560 17248 7560 17248 0 _1350_
rlabel via2 17304 18312 17304 18312 0 _1351_
rlabel metal2 17864 19880 17864 19880 0 _1352_
rlabel metal2 7280 16856 7280 16856 0 _1353_
rlabel metal2 7112 26264 7112 26264 0 _1354_
rlabel metal2 11592 8960 11592 8960 0 _1355_
rlabel metal2 10696 7224 10696 7224 0 _1356_
rlabel metal2 11872 2856 11872 2856 0 _1357_
rlabel metal2 11984 11368 11984 11368 0 _1358_
rlabel metal2 15960 8288 15960 8288 0 _1359_
rlabel metal2 16240 9240 16240 9240 0 _1360_
rlabel metal3 20048 10584 20048 10584 0 _1361_
rlabel metal2 15288 20104 15288 20104 0 _1362_
rlabel metal2 20832 22232 20832 22232 0 _1363_
rlabel metal3 26096 15176 26096 15176 0 _1364_
rlabel metal2 7840 24584 7840 24584 0 _1365_
rlabel metal2 10024 20272 10024 20272 0 _1366_
rlabel metal2 22624 18424 22624 18424 0 _1367_
rlabel metal2 19264 25368 19264 25368 0 _1368_
rlabel metal2 6888 18872 6888 18872 0 _1369_
rlabel metal2 27608 15680 27608 15680 0 _1370_
rlabel metal2 27328 21896 27328 21896 0 _1371_
rlabel metal2 29176 21280 29176 21280 0 _1372_
rlabel metal2 26600 20048 26600 20048 0 _1373_
rlabel metal2 17976 16912 17976 16912 0 _1374_
rlabel metal2 17752 17192 17752 17192 0 _1375_
rlabel metal2 18200 22512 18200 22512 0 _1376_
rlabel metal2 26936 16800 26936 16800 0 _1377_
rlabel metal2 23128 23184 23128 23184 0 _1378_
rlabel metal3 13328 25480 13328 25480 0 _1379_
rlabel metal2 17080 21840 17080 21840 0 _1380_
rlabel metal2 24024 20608 24024 20608 0 _1381_
rlabel metal2 29848 21560 29848 21560 0 _1382_
rlabel metal2 27944 20776 27944 20776 0 _1383_
rlabel metal3 25256 20104 25256 20104 0 _1384_
rlabel metal2 33656 19936 33656 19936 0 _1385_
rlabel metal2 42000 23128 42000 23128 0 _1386_
rlabel metal2 15512 17976 15512 17976 0 _1387_
rlabel metal3 44016 23688 44016 23688 0 _1388_
rlabel metal3 35280 22344 35280 22344 0 _1389_
rlabel metal2 45416 23072 45416 23072 0 _1390_
rlabel metal2 45528 22512 45528 22512 0 _1391_
rlabel metal2 45976 23688 45976 23688 0 _1392_
rlabel metal2 46648 24416 46648 24416 0 _1393_
rlabel metal2 46872 25144 46872 25144 0 _1394_
rlabel metal2 47264 24136 47264 24136 0 _1395_
rlabel metal3 48496 23128 48496 23128 0 _1396_
rlabel metal2 31304 25648 31304 25648 0 _1397_
rlabel metal2 30968 21504 30968 21504 0 _1398_
rlabel metal3 16912 27048 16912 27048 0 _1399_
rlabel metal2 19488 23352 19488 23352 0 _1400_
rlabel metal2 14168 22736 14168 22736 0 _1401_
rlabel metal2 12040 19656 12040 19656 0 _1402_
rlabel metal3 22400 15848 22400 15848 0 _1403_
rlabel metal2 21784 25928 21784 25928 0 _1404_
rlabel metal2 32088 24416 32088 24416 0 _1405_
rlabel metal3 24976 22344 24976 22344 0 _1406_
rlabel metal2 18984 18536 18984 18536 0 _1407_
rlabel metal2 27664 23912 27664 23912 0 _1408_
rlabel metal2 18984 20720 18984 20720 0 _1409_
rlabel metal2 29960 22848 29960 22848 0 _1410_
rlabel metal2 31416 22512 31416 22512 0 _1411_
rlabel metal2 43512 24136 43512 24136 0 _1412_
rlabel metal3 44632 23240 44632 23240 0 _1413_
rlabel metal2 35112 24584 35112 24584 0 _1414_
rlabel metal2 18704 20552 18704 20552 0 _1415_
rlabel metal2 19208 4816 19208 4816 0 _1416_
rlabel metal2 14840 22736 14840 22736 0 _1417_
rlabel metal2 15736 23856 15736 23856 0 _1418_
rlabel metal2 29344 24920 29344 24920 0 _1419_
rlabel metal2 26936 22848 26936 22848 0 _1420_
rlabel metal2 26376 23576 26376 23576 0 _1421_
rlabel metal2 21672 20496 21672 20496 0 _1422_
rlabel metal3 24080 23016 24080 23016 0 _1423_
rlabel metal2 26096 23240 26096 23240 0 _1424_
rlabel metal2 31976 22736 31976 22736 0 _1425_
rlabel metal3 33096 23128 33096 23128 0 _1426_
rlabel metal2 37016 22904 37016 22904 0 _1427_
rlabel metal2 33824 16856 33824 16856 0 _1428_
rlabel metal2 25872 24024 25872 24024 0 _1429_
rlabel metal3 7784 23912 7784 23912 0 _1430_
rlabel metal3 25200 21784 25200 21784 0 _1431_
rlabel metal2 27272 17360 27272 17360 0 _1432_
rlabel metal2 18200 17304 18200 17304 0 _1433_
rlabel metal2 14728 17640 14728 17640 0 _1434_
rlabel metal3 19208 1400 19208 1400 0 _1435_
rlabel metal3 20328 21616 20328 21616 0 _1436_
rlabel metal2 20216 21896 20216 21896 0 _1437_
rlabel metal2 15512 24976 15512 24976 0 _1438_
rlabel metal2 16296 20552 16296 20552 0 _1439_
rlabel metal2 21112 21616 21112 21616 0 _1440_
rlabel metal2 10808 19040 10808 19040 0 _1441_
rlabel metal2 1960 27440 1960 27440 0 addI[0]
rlabel metal3 1358 28280 1358 28280 0 addI[1]
rlabel metal3 1638 29624 1638 29624 0 addI[2]
rlabel metal3 1358 28952 1358 28952 0 addI[3]
rlabel metal3 1358 30296 1358 30296 0 addI[4]
rlabel metal3 29512 3416 29512 3416 0 addI[5]
rlabel metal3 1358 35000 1358 35000 0 addQ[0]
rlabel metal3 1358 36344 1358 36344 0 addQ[1]
rlabel metal3 1358 47768 1358 47768 0 addQ[2]
rlabel metal3 1358 48440 1358 48440 0 addQ[3]
rlabel metal3 1358 54488 1358 54488 0 addQ[4]
rlabel metal2 30968 57610 30968 57610 0 addQ[5]
rlabel metal3 32536 29624 32536 29624 0 bit2symb.regi
rlabel metal3 19320 31080 19320 31080 0 clknet_0_CLK
rlabel metal3 16408 33320 16408 33320 0 clknet_1_0__leaf_CLK
rlabel metal2 25032 30968 25032 30968 0 clknet_1_1__leaf_CLK
rlabel metal2 33992 30632 33992 30632 0 net1
rlabel metal2 53032 18312 53032 18312 0 net10
rlabel metal3 1470 25592 1470 25592 0 net100
rlabel metal3 1246 42392 1246 42392 0 net101
rlabel metal2 58184 10640 58184 10640 0 net102
rlabel metal2 8792 57610 8792 57610 0 net103
rlabel metal3 1470 37016 1470 37016 0 net104
rlabel metal2 53032 16016 53032 16016 0 net11
rlabel metal2 53368 14952 53368 14952 0 net12
rlabel metal2 51688 11312 51688 11312 0 net13
rlabel metal2 52024 8176 52024 8176 0 net14
rlabel metal2 51072 5992 51072 5992 0 net15
rlabel metal3 51128 4872 51128 4872 0 net16
rlabel metal3 42168 56056 42168 56056 0 net17
rlabel metal2 55608 35392 55608 35392 0 net18
rlabel metal2 54376 33264 54376 33264 0 net19
rlabel metal2 17528 31360 17528 31360 0 net2
rlabel metal2 55832 36736 55832 36736 0 net20
rlabel metal3 46984 56056 46984 56056 0 net21
rlabel metal3 53536 56056 53536 56056 0 net22
rlabel metal2 53928 53648 53928 53648 0 net23
rlabel metal2 55272 49056 55272 49056 0 net24
rlabel metal2 55272 50512 55272 50512 0 net25
rlabel metal2 55944 44744 55944 44744 0 net26
rlabel metal2 56056 43176 56056 43176 0 net27
rlabel metal2 56056 40824 56056 40824 0 net28
rlabel metal2 56056 38528 56056 38528 0 net29
rlabel metal2 7560 34776 7560 34776 0 net3
rlabel metal2 7784 29344 7784 29344 0 net30
rlabel metal2 7336 27328 7336 27328 0 net31
rlabel metal2 8456 29624 8456 29624 0 net32
rlabel metal3 15624 29344 15624 29344 0 net33
rlabel metal2 21336 31192 21336 31192 0 net34
rlabel metal2 29064 3584 29064 3584 0 net35
rlabel metal2 9464 35896 9464 35896 0 net36
rlabel metal2 9744 36456 9744 36456 0 net37
rlabel metal2 4312 47768 4312 47768 0 net38
rlabel metal3 5208 48776 5208 48776 0 net39
rlabel metal2 47096 25424 47096 25424 0 net4
rlabel metal2 4200 55160 4200 55160 0 net40
rlabel metal3 30800 32760 30800 32760 0 net41
rlabel metal2 39816 28504 39816 28504 0 net42
rlabel metal2 39256 26320 39256 26320 0 net43
rlabel metal2 39760 26488 39760 26488 0 net44
rlabel metal2 27496 6384 27496 6384 0 net45
rlabel metal4 25704 40208 25704 40208 0 net46
rlabel metal2 40936 33432 40936 33432 0 net47
rlabel metal2 42728 30184 42728 30184 0 net48
rlabel metal2 23576 53424 23576 53424 0 net49
rlabel metal2 47488 4872 47488 4872 0 net5
rlabel metal2 8008 39424 8008 39424 0 net50
rlabel metal3 5768 37240 5768 37240 0 net51
rlabel metal2 10136 35616 10136 35616 0 net52
rlabel metal2 16408 28672 16408 28672 0 net53
rlabel metal2 8120 25872 8120 25872 0 net54
rlabel metal2 4872 26572 4872 26572 0 net55
rlabel metal2 8344 34496 8344 34496 0 net56
rlabel metal2 9128 31472 9128 31472 0 net57
rlabel metal3 8960 34776 8960 34776 0 net58
rlabel metal2 22008 31640 22008 31640 0 net59
rlabel metal2 43624 4368 43624 4368 0 net6
rlabel metal2 30856 29792 30856 29792 0 net60
rlabel metal3 44800 28056 44800 28056 0 net61
rlabel metal3 43680 31192 43680 31192 0 net62
rlabel metal2 37352 29792 37352 29792 0 net63
rlabel metal2 43456 33096 43456 33096 0 net64
rlabel metal2 43176 32872 43176 32872 0 net65
rlabel metal2 10920 33712 10920 33712 0 net66
rlabel metal2 58184 47152 58184 47152 0 net67
rlabel metal2 58184 13664 58184 13664 0 net68
rlabel metal2 7560 56280 7560 56280 0 net69
rlabel metal2 43848 5096 43848 5096 0 net7
rlabel metal2 58184 28336 58184 28336 0 net70
rlabel metal2 57736 10416 57736 10416 0 net71
rlabel metal2 6216 56280 6216 56280 0 net72
rlabel metal3 1246 39032 1246 39032 0 net73
rlabel metal2 58184 18928 58184 18928 0 net74
rlabel metal3 1246 17528 1246 17528 0 net75
rlabel metal2 10920 56280 10920 56280 0 net76
rlabel metal3 1246 51128 1246 51128 0 net77
rlabel metal2 58240 26824 58240 26824 0 net78
rlabel metal2 58184 25984 58184 25984 0 net79
rlabel metal2 50120 23856 50120 23856 0 net8
rlabel metal3 1246 35672 1246 35672 0 net80
rlabel metal3 1582 31640 1582 31640 0 net81
rlabel metal2 58184 9520 58184 9520 0 net82
rlabel metal2 58184 16576 58184 16576 0 net83
rlabel metal2 58184 22008 58184 22008 0 net84
rlabel metal2 55048 56448 55048 56448 0 net85
rlabel metal2 9464 2030 9464 2030 0 net86
rlabel metal3 1246 20888 1246 20888 0 net87
rlabel metal2 9576 56280 9576 56280 0 net88
rlabel metal2 58184 7896 58184 7896 0 net89
rlabel metal2 51128 22064 51128 22064 0 net9
rlabel metal2 52472 2030 52472 2030 0 net90
rlabel metal3 58744 20216 58744 20216 0 net91
rlabel metal2 55160 57778 55160 57778 0 net92
rlabel metal2 4760 2030 4760 2030 0 net93
rlabel metal2 1736 26712 1736 26712 0 net94
rlabel metal2 58184 12432 58184 12432 0 net95
rlabel metal2 11592 56280 11592 56280 0 net96
rlabel metal2 5544 56280 5544 56280 0 net97
rlabel metal3 1246 24248 1246 24248 0 net98
rlabel metal3 1246 41048 1246 41048 0 net99
rlabel metal3 42336 24808 42336 24808 0 p_shaping_I.bit_in
rlabel metal2 32368 21672 32368 21672 0 p_shaping_I.bit_in_1
rlabel metal2 34440 26152 34440 26152 0 p_shaping_I.bit_in_2
rlabel metal2 43512 25312 43512 25312 0 p_shaping_I.counter\[0\]
rlabel metal2 41776 23912 41776 23912 0 p_shaping_I.counter\[1\]
rlabel metal2 38416 27944 38416 27944 0 p_shaping_I.ctl_1
rlabel metal2 41944 47768 41944 47768 0 p_shaping_Q.bit_in_1
rlabel metal2 44016 48104 44016 48104 0 p_shaping_Q.bit_in_2
rlabel metal2 45976 30576 45976 30576 0 p_shaping_Q.counter\[0\]
rlabel metal3 46536 48104 46536 48104 0 p_shaping_Q.counter\[1\]
rlabel metal2 42168 30688 42168 30688 0 p_shaping_Q.ctl_1
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
