VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO OQPSK_PS_RCOSINE2
  CLASS BLOCK ;
  FOREIGN OQPSK_PS_RCOSINE2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN BitIn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 151.200 300.000 151.760 ;
    END
  END BitIn
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 168.000 4.000 168.560 ;
    END
  END CLK
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 154.560 4.000 155.120 ;
    END
  END EN
  PIN I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 124.320 300.000 124.880 ;
    END
  END I[0]
  PIN I[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 231.840 0.000 232.400 4.000 ;
    END
  END I[10]
  PIN I[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 0.000 218.960 4.000 ;
    END
  END I[11]
  PIN I[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 211.680 0.000 212.240 4.000 ;
    END
  END I[12]
  PIN I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 117.600 300.000 118.160 ;
    END
  END I[1]
  PIN I[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 107.520 300.000 108.080 ;
    END
  END I[2]
  PIN I[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 90.720 300.000 91.280 ;
    END
  END I[3]
  PIN I[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 84.000 300.000 84.560 ;
    END
  END I[4]
  PIN I[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 77.280 300.000 77.840 ;
    END
  END I[5]
  PIN I[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 57.120 300.000 57.680 ;
    END
  END I[6]
  PIN I[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 43.680 300.000 44.240 ;
    END
  END I[7]
  PIN I[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 255.360 0.000 255.920 4.000 ;
    END
  END I[8]
  PIN I[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 252.000 0.000 252.560 4.000 ;
    END
  END I[9]
  PIN Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 296.000 205.520 300.000 ;
    END
  END Q[0]
  PIN Q[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 174.720 300.000 175.280 ;
    END
  END Q[10]
  PIN Q[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 164.640 300.000 165.200 ;
    END
  END Q[11]
  PIN Q[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 178.080 300.000 178.640 ;
    END
  END Q[12]
  PIN Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 228.480 296.000 229.040 300.000 ;
    END
  END Q[1]
  PIN Q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 296.000 262.640 300.000 ;
    END
  END Q[2]
  PIN Q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 265.440 300.000 266.000 ;
    END
  END Q[3]
  PIN Q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 252.000 300.000 252.560 ;
    END
  END Q[4]
  PIN Q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 248.640 300.000 249.200 ;
    END
  END Q[5]
  PIN Q[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 221.760 300.000 222.320 ;
    END
  END Q[6]
  PIN Q[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 215.040 300.000 215.600 ;
    END
  END Q[7]
  PIN Q[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 201.600 300.000 202.160 ;
    END
  END Q[8]
  PIN Q[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 188.160 300.000 188.720 ;
    END
  END Q[9]
  PIN RST
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 164.640 4.000 165.200 ;
    END
  END RST
  PIN addI[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 137.760 4.000 138.320 ;
    END
  END addI[0]
  PIN addI[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 141.120 4.000 141.680 ;
    END
  END addI[1]
  PIN addI[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 147.840 4.000 148.400 ;
    END
  END addI[2]
  PIN addI[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 144.480 4.000 145.040 ;
    END
  END addI[3]
  PIN addI[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 151.200 4.000 151.760 ;
    END
  END addI[4]
  PIN addI[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 0.000 145.040 4.000 ;
    END
  END addI[5]
  PIN addQ[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 174.720 4.000 175.280 ;
    END
  END addQ[0]
  PIN addQ[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 181.440 4.000 182.000 ;
    END
  END addQ[1]
  PIN addQ[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 238.560 4.000 239.120 ;
    END
  END addQ[2]
  PIN addQ[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 241.920 4.000 242.480 ;
    END
  END addQ[3]
  PIN addQ[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 272.160 4.000 272.720 ;
    END
  END addQ[4]
  PIN addQ[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 296.000 155.120 300.000 ;
    END
  END addQ[5]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 120.960 4.000 121.520 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 141.120 300.000 141.680 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 50.400 300.000 50.960 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 296.000 30.800 300.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 194.880 4.000 195.440 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 94.080 300.000 94.640 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 87.360 4.000 87.920 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 296.000 54.320 300.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 255.360 4.000 255.920 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 131.040 300.000 131.600 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 127.680 300.000 128.240 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 204.960 4.000 205.520 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 178.080 4.000 178.640 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 157.920 4.000 158.480 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 47.040 300.000 47.600 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 80.640 300.000 81.200 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 110.880 300.000 111.440 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 272.160 296.000 272.720 300.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 0.000 47.600 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 104.160 4.000 104.720 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 296.000 47.600 300.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 40.320 300.000 40.880 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 127.680 4.000 128.240 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 0.000 262.640 4.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 97.440 300.000 98.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 275.520 296.000 276.080 300.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 0.000 24.080 4.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 134.400 4.000 134.960 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 60.480 300.000 61.040 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 296.000 57.680 300.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 296.000 27.440 300.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 211.680 4.000 212.240 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 53.760 300.000 54.320 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 296.000 44.240 300.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 184.800 4.000 185.360 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 235.200 300.000 235.760 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 67.200 300.000 67.760 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 296.000 37.520 300.000 ;
    END
  END io_oeb[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 282.540 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 282.540 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 292.880 283.210 ;
      LAYER Metal2 ;
        RECT 8.540 295.700 26.580 296.000 ;
        RECT 27.740 295.700 29.940 296.000 ;
        RECT 31.100 295.700 36.660 296.000 ;
        RECT 37.820 295.700 43.380 296.000 ;
        RECT 44.540 295.700 46.740 296.000 ;
        RECT 47.900 295.700 53.460 296.000 ;
        RECT 54.620 295.700 56.820 296.000 ;
        RECT 57.980 295.700 154.260 296.000 ;
        RECT 155.420 295.700 204.660 296.000 ;
        RECT 205.820 295.700 228.180 296.000 ;
        RECT 229.340 295.700 261.780 296.000 ;
        RECT 262.940 295.700 271.860 296.000 ;
        RECT 273.020 295.700 275.220 296.000 ;
        RECT 276.380 295.700 291.620 296.000 ;
        RECT 8.540 4.300 291.620 295.700 ;
        RECT 8.540 4.000 23.220 4.300 ;
        RECT 24.380 4.000 46.740 4.300 ;
        RECT 47.900 4.000 144.180 4.300 ;
        RECT 145.340 4.000 211.380 4.300 ;
        RECT 212.540 4.000 218.100 4.300 ;
        RECT 219.260 4.000 231.540 4.300 ;
        RECT 232.700 4.000 251.700 4.300 ;
        RECT 252.860 4.000 255.060 4.300 ;
        RECT 256.220 4.000 261.780 4.300 ;
        RECT 262.940 4.000 291.620 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 273.020 296.660 289.380 ;
        RECT 4.300 271.860 296.660 273.020 ;
        RECT 4.000 266.300 296.660 271.860 ;
        RECT 4.000 265.140 295.700 266.300 ;
        RECT 4.000 256.220 296.660 265.140 ;
        RECT 4.300 255.060 296.660 256.220 ;
        RECT 4.000 252.860 296.660 255.060 ;
        RECT 4.000 251.700 295.700 252.860 ;
        RECT 4.000 249.500 296.660 251.700 ;
        RECT 4.000 248.340 295.700 249.500 ;
        RECT 4.000 242.780 296.660 248.340 ;
        RECT 4.300 241.620 296.660 242.780 ;
        RECT 4.000 239.420 296.660 241.620 ;
        RECT 4.300 238.260 296.660 239.420 ;
        RECT 4.000 236.060 296.660 238.260 ;
        RECT 4.000 234.900 295.700 236.060 ;
        RECT 4.000 222.620 296.660 234.900 ;
        RECT 4.000 221.460 295.700 222.620 ;
        RECT 4.000 215.900 296.660 221.460 ;
        RECT 4.000 214.740 295.700 215.900 ;
        RECT 4.000 212.540 296.660 214.740 ;
        RECT 4.300 211.380 296.660 212.540 ;
        RECT 4.000 205.820 296.660 211.380 ;
        RECT 4.300 204.660 296.660 205.820 ;
        RECT 4.000 202.460 296.660 204.660 ;
        RECT 4.000 201.300 295.700 202.460 ;
        RECT 4.000 195.740 296.660 201.300 ;
        RECT 4.300 194.580 296.660 195.740 ;
        RECT 4.000 189.020 296.660 194.580 ;
        RECT 4.000 187.860 295.700 189.020 ;
        RECT 4.000 185.660 296.660 187.860 ;
        RECT 4.300 184.500 296.660 185.660 ;
        RECT 4.000 182.300 296.660 184.500 ;
        RECT 4.300 181.140 296.660 182.300 ;
        RECT 4.000 178.940 296.660 181.140 ;
        RECT 4.300 177.780 295.700 178.940 ;
        RECT 4.000 175.580 296.660 177.780 ;
        RECT 4.300 174.420 295.700 175.580 ;
        RECT 4.000 168.860 296.660 174.420 ;
        RECT 4.300 167.700 296.660 168.860 ;
        RECT 4.000 165.500 296.660 167.700 ;
        RECT 4.300 164.340 295.700 165.500 ;
        RECT 4.000 158.780 296.660 164.340 ;
        RECT 4.300 157.620 296.660 158.780 ;
        RECT 4.000 155.420 296.660 157.620 ;
        RECT 4.300 154.260 296.660 155.420 ;
        RECT 4.000 152.060 296.660 154.260 ;
        RECT 4.300 150.900 295.700 152.060 ;
        RECT 4.000 148.700 296.660 150.900 ;
        RECT 4.300 147.540 296.660 148.700 ;
        RECT 4.000 145.340 296.660 147.540 ;
        RECT 4.300 144.180 296.660 145.340 ;
        RECT 4.000 141.980 296.660 144.180 ;
        RECT 4.300 140.820 295.700 141.980 ;
        RECT 4.000 138.620 296.660 140.820 ;
        RECT 4.300 137.460 296.660 138.620 ;
        RECT 4.000 135.260 296.660 137.460 ;
        RECT 4.300 134.100 296.660 135.260 ;
        RECT 4.000 131.900 296.660 134.100 ;
        RECT 4.000 130.740 295.700 131.900 ;
        RECT 4.000 128.540 296.660 130.740 ;
        RECT 4.300 127.380 295.700 128.540 ;
        RECT 4.000 125.180 296.660 127.380 ;
        RECT 4.000 124.020 295.700 125.180 ;
        RECT 4.000 121.820 296.660 124.020 ;
        RECT 4.300 120.660 296.660 121.820 ;
        RECT 4.000 118.460 296.660 120.660 ;
        RECT 4.000 117.300 295.700 118.460 ;
        RECT 4.000 111.740 296.660 117.300 ;
        RECT 4.000 110.580 295.700 111.740 ;
        RECT 4.000 108.380 296.660 110.580 ;
        RECT 4.000 107.220 295.700 108.380 ;
        RECT 4.000 105.020 296.660 107.220 ;
        RECT 4.300 103.860 296.660 105.020 ;
        RECT 4.000 98.300 296.660 103.860 ;
        RECT 4.000 97.140 295.700 98.300 ;
        RECT 4.000 94.940 296.660 97.140 ;
        RECT 4.000 93.780 295.700 94.940 ;
        RECT 4.000 91.580 296.660 93.780 ;
        RECT 4.000 90.420 295.700 91.580 ;
        RECT 4.000 88.220 296.660 90.420 ;
        RECT 4.300 87.060 296.660 88.220 ;
        RECT 4.000 84.860 296.660 87.060 ;
        RECT 4.000 83.700 295.700 84.860 ;
        RECT 4.000 81.500 296.660 83.700 ;
        RECT 4.000 80.340 295.700 81.500 ;
        RECT 4.000 78.140 296.660 80.340 ;
        RECT 4.000 76.980 295.700 78.140 ;
        RECT 4.000 68.060 296.660 76.980 ;
        RECT 4.000 66.900 295.700 68.060 ;
        RECT 4.000 61.340 296.660 66.900 ;
        RECT 4.000 60.180 295.700 61.340 ;
        RECT 4.000 57.980 296.660 60.180 ;
        RECT 4.000 56.820 295.700 57.980 ;
        RECT 4.000 54.620 296.660 56.820 ;
        RECT 4.000 53.460 295.700 54.620 ;
        RECT 4.000 51.260 296.660 53.460 ;
        RECT 4.000 50.100 295.700 51.260 ;
        RECT 4.000 47.900 296.660 50.100 ;
        RECT 4.000 46.740 295.700 47.900 ;
        RECT 4.000 44.540 296.660 46.740 ;
        RECT 4.000 43.380 295.700 44.540 ;
        RECT 4.000 41.180 296.660 43.380 ;
        RECT 4.000 40.020 295.700 41.180 ;
        RECT 4.000 6.860 296.660 40.020 ;
      LAYER Metal4 ;
        RECT 34.300 282.840 232.820 289.430 ;
        RECT 34.300 15.080 98.740 282.840 ;
        RECT 100.940 15.080 175.540 282.840 ;
        RECT 177.740 15.080 232.820 282.840 ;
        RECT 34.300 6.810 232.820 15.080 ;
  END
END OQPSK_PS_RCOSINE2
END LIBRARY

