// This is the unpowered netlist.
module OQPSK_PS_RCOSINE2 (BitIn,
    CLK,
    EN,
    RST,
    I,
    Q,
    addI,
    addQ,
    io_oeb);
 input BitIn;
 input CLK;
 input EN;
 input RST;
 output [12:0] I;
 output [12:0] Q;
 output [5:0] addI;
 output [5:0] addQ;
 output [37:0] io_oeb;

 wire net98;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net99;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net100;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net67;
 wire net68;
 wire net69;
 wire \Reg_Delay_Q.In ;
 wire \Reg_Delay_Q.Out ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire \bit2symb.regi ;
 wire clknet_0_CLK;
 wire clknet_1_0__leaf_CLK;
 wire clknet_1_1__leaf_CLK;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net7;
 wire net8;
 wire net9;
 wire \p_shaping_I.bit_in ;
 wire \p_shaping_I.bit_in_1 ;
 wire \p_shaping_I.bit_in_2 ;
 wire \p_shaping_I.counter[0] ;
 wire \p_shaping_I.counter[1] ;
 wire \p_shaping_I.ctl_1 ;
 wire \p_shaping_Q.bit_in_1 ;
 wire \p_shaping_Q.bit_in_2 ;
 wire \p_shaping_Q.counter[0] ;
 wire \p_shaping_Q.counter[1] ;
 wire \p_shaping_Q.ctl_1 ;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1455__A1 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1456__I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1457__A1 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1468__I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1469__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1470__A1 (.I(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1474__A2 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1475__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1477__A1 (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1478__A2 (.I(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1478__B (.I(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1478__C (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1479__A1 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1487__I (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1488__I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1494__A1 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1497__I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1500__I (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1504__A1 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1504__A2 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1506__I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1508__A2 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1509__B (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1513__I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1520__A1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1520__A2 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1520__B (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1521__A1 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1521__A3 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1523__I (.I(\p_shaping_I.bit_in_1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1531__A1 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1534__I (.I(\p_shaping_Q.bit_in_1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1545__I (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1558__I (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1559__A2 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1564__I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1567__I (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1571__A1 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1571__B (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1575__B2 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1581__I (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1584__I (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1587__A2 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1587__B (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1588__A2 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1588__B (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1589__A1 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1590__A1 (.I(\p_shaping_Q.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1591__I (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1594__I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1595__I (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1601__A2 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1605__A1 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1606__A2 (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1607__A3 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1607__B (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1611__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1611__B (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1612__I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1615__A3 (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1617__A1 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1618__A1 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1619__I0 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1620__I (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1622__I (.I(\p_shaping_Q.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1625__I (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1627__I (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1636__A2 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1642__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1642__B (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1643__A1 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1645__A1 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1645__B1 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1646__A1 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1646__A2 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1648__A1 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1649__A1 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1654__I (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1655__I (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1656__I (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1657__I (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1658__A3 (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1659__A2 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1660__A2 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1660__B1 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1663__A1 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1663__B (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1665__I (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1666__A2 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1667__A1 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1669__A1 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1669__A2 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1672__A1 (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1672__C2 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1673__A1 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1675__A1 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1676__I (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1678__A2 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1679__A1 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1683__A1 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1688__I1 (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1688__S0 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1690__A1 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1693__I (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1695__A1 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1695__A2 (.I(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1695__B (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1697__A1 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1698__C (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1701__A2 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1702__B (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1705__A1 (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1705__C (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1706__A2 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1707__A1 (.I(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1710__I (.I(\p_shaping_Q.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1714__B (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1718__A3 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1721__A1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1721__A2 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1722__A1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1722__A2 (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1723__A1 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1725__A2 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1725__A3 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1727__I (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1728__I (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1735__I (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1736__A2 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1736__A3 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1737__A2 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1741__A1 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1743__B (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1746__A1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1746__A2 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1747__A2 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1749__A2 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1749__B (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1761__A1 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1763__A1 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1765__A2 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1766__I (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1767__A1 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1772__A2 (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1775__A2 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1779__A1 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1784__I (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1785__I (.I(\p_shaping_Q.bit_in_1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1786__C (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1793__A1 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1793__A2 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1795__A1 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1796__A2 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1796__B (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1797__A1 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1798__B (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1799__A2 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1800__A1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1805__A1 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1805__A2 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1808__A2 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1813__A1 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1818__B1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1820__A1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1831__B (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1835__A2 (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1837__A1 (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1837__A2 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1838__A2 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1839__A1 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1840__A1 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1841__B2 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1843__A2 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1843__B (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1844__B (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1852__A1 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1852__A2 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1854__A2 (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1855__A2 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1857__A3 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1860__C (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1862__B2 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1864__A1 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1866__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1870__A1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1870__A2 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1871__A1 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1872__A2 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1873__C (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1874__A1 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1874__A3 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1879__A1 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1883__I (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1884__A1 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1892__A1 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1892__A2 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1897__B2 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1897__C (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1898__I (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1899__I (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1901__A1 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1907__A1 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1910__A3 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1911__A1 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1914__A1 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1917__A1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1918__I (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1921__A1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1921__A4 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1923__B (.I(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1925__A2 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1927__A1 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1928__A2 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1931__A1 (.I(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1932__A2 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1946__A1 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1950__I (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1951__A3 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1952__B (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1955__A1 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1959__A3 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1959__A4 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1960__A2 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1960__B (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1963__A2 (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1965__A1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1970__A1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1970__A4 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1972__A2 (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1975__A2 (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1975__A3 (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1976__A1 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1976__A2 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1977__A2 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1977__B (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1978__A1 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1978__A3 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1979__A1 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1980__C (.I(\p_shaping_Q.bit_in_1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1983__A1 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2001__I (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2002__B (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2006__A2 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2007__A1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2007__A2 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2012__A1 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2013__A2 (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2017__A2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2018__A1 (.I(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2018__B2 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2019__A2 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2021__A1 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2021__A2 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2022__A1 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2022__A2 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2024__A1 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2026__A2 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2034__A2 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2036__S (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2037__B (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2051__A1 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2062__A1 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2062__B1 (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2065__A1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2067__A1 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2074__C (.I(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2080__A1 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2080__B (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2096__A1 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2097__A1 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2099__A2 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2100__B2 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2101__A1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2102__A3 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2108__A1 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2111__A2 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2112__A1 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2117__A2 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2119__B (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2129__A1 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2132__A1 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2134__B (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2137__A2 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2138__A2 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2139__A2 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2164__A2 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2171__I (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2187__A2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2190__A1 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2190__C (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2207__B2 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2216__B (.I(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2223__I (.I(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2228__A2 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2234__A1 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2234__A2 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2234__C1 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2238__I (.I(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2244__B (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2249__C (.I(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2255__A2 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2258__B (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2261__A2 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2269__A1 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2269__B1 (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2270__A1 (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2289__A2 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2289__B (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2291__I (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2292__I (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2294__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2294__A3 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2297__A1 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2297__A2 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2299__I (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2300__A2 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2300__A3 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2303__A2 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2313__I (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2322__A1 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2322__A2 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2327__I0 (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2327__I3 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2327__S1 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2330__A1 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2331__A1 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2331__A2 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2335__A2 (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2339__A2 (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2339__B1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2339__B2 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2341__A1 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2343__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2343__A2 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2350__A2 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2359__A2 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2362__A3 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2366__A1 (.I(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2367__A2 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2369__A2 (.I(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2370__A2 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2371__A3 (.I(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2373__A1 (.I(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2375__A2 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2378__A2 (.I(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2381__A2 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2382__A2 (.I(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2382__A3 (.I(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2384__I (.I(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2385__A2 (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2387__I (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__C (.I(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2392__A4 (.I(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2393__I (.I(\p_shaping_I.bit_in_1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2395__A1 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2397__B (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2398__A3 (.I(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2404__A2 (.I(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2405__A2 (.I(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2405__A3 (.I(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2407__A1 (.I(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2409__A1 (.I(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2413__B2 (.I(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2427__A1 (.I(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2430__A1 (.I(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2430__A2 (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2431__A1 (.I(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2436__I (.I(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2437__A1 (.I(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2437__B (.I(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__A2 (.I(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2444__A1 (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2444__B1 (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2444__B2 (.I(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__A1 (.I(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__A2 (.I(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2446__C (.I(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2448__B (.I(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2449__A3 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2450__A2 (.I(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2451__A1 (.I(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2451__A2 (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2453__A2 (.I(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2454__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2454__A2 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2456__A2 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2457__A2 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2459__A1 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2459__B (.I(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2460__A1 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2461__A1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2461__A2 (.I(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2462__A3 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2463__A1 (.I(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2464__I (.I(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__A2 (.I(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2468__A2 (.I(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2473__A3 (.I(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2476__I0 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2476__S (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2477__A2 (.I(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2478__A1 (.I(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2487__A2 (.I(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2497__I (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2499__A2 (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2500__A1 (.I(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2501__I (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2502__A1 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2502__B (.I(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2503__A2 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2504__B1 (.I(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2504__B2 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2507__A2 (.I(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2508__A1 (.I(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2508__B2 (.I(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2510__A2 (.I(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2511__A1 (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__C (.I(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__A1 (.I(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__A1 (.I(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__A2 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2519__A1 (.I(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__A2 (.I(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__B (.I(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__A1 (.I(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2525__A1 (.I(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2525__B (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2526__A2 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2527__B (.I(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2528__A1 (.I(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2529__A1 (.I(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2530__A3 (.I(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2532__A3 (.I(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2533__A1 (.I(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__A2 (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2537__A2 (.I(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2540__A3 (.I(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2547__A1 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2549__I (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2551__A1 (.I(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2561__A2 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2561__B (.I(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2562__A1 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2562__A2 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2564__A2 (.I(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2565__A2 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2566__A1 (.I(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2567__C (.I(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2568__A1 (.I(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2569__A2 (.I(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2569__A3 (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2571__A1 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2572__A1 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2575__B (.I(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2575__C (.I(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__A2 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2577__A1 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2585__A1 (.I(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2586__B (.I(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2588__A2 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2588__B (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2589__A1 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2589__A3 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2597__I (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2598__I (.I(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2600__A1 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2600__B (.I(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2601__I (.I(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2602__A1 (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2604__A2 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2609__A2 (.I(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2610__A2 (.I(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2611__A1 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2611__B2 (.I(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2631__A2 (.I(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2631__A3 (.I(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2635__I (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__A2 (.I(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__A1 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__A2 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2640__A1 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2642__A1 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2644__A1 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2644__A2 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2645__A2 (.I(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2646__A2 (.I(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2649__A1 (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2649__C (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2667__B (.I(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2676__A1 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2680__A1 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2680__A2 (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2680__C (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2682__I (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2689__I (.I(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2691__A2 (.I(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2692__A1 (.I(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2692__A2 (.I(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2693__A2 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2693__B2 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2694__A1 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2696__A1 (.I(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2699__A2 (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2699__A3 (.I(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2700__A2 (.I(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2701__A1 (.I(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2702__A3 (.I(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2703__A2 (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2706__A2 (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2722__A1 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2722__A2 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2723__A2 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2724__A2 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2725__A3 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2731__A2 (.I(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2732__B (.I(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2733__B (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2734__B2 (.I(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2735__A2 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2736__A2 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2742__A2 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__A2 (.I(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2745__A1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2745__A2 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2746__A1 (.I(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2760__A2 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2760__A3 (.I(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2762__B (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2765__A1 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2767__A1 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2773__A1 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2776__S (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2788__A1 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2788__A2 (.I(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2789__A1 (.I(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2789__A2 (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2790__I0 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2791__I (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2792__A2 (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2793__B (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2794__A1 (.I(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2794__A2 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2794__C (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__A1 (.I(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__A2 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__B (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2799__A1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2803__C (.I(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2817__A1 (.I(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2818__A2 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2822__A2 (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2823__A1 (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2823__C (.I(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2837__A1 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2837__B (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2863__A1 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2864__I1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2866__A1 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2867__I (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2871__A1 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2874__A2 (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2875__A1 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2875__B1 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2876__A2 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2880__A1 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2882__A1 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2883__A1 (.I(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2883__A2 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2884__A1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2885__A2 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2888__A2 (.I(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2888__B2 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2889__A1 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2892__A1 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2893__A1 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2894__A1 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2894__B1 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2895__A1 (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2895__A2 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2897__A2 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2897__A3 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2900__A1 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2900__A2 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2902__A2 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2906__I1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2908__A1 (.I(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2909__A1 (.I(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2913__CLK (.I(clknet_1_0__leaf_CLK));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2914__CLK (.I(clknet_1_0__leaf_CLK));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2915__CLK (.I(clknet_1_0__leaf_CLK));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2916__CLK (.I(clknet_1_0__leaf_CLK));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2919__CLK (.I(clknet_1_0__leaf_CLK));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2920__CLK (.I(clknet_1_0__leaf_CLK));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2921__CLK (.I(clknet_1_0__leaf_CLK));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2922__CLK (.I(clknet_1_0__leaf_CLK));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2923__CLK (.I(clknet_1_0__leaf_CLK));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2929__D (.I(\p_shaping_I.bit_in_1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2929__RN (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2933__D (.I(\p_shaping_Q.bit_in_1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2935__D (.I(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_CLK_I (.I(CLK));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout42_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout43_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout49_I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout50_I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout59_I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout60_I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout63_I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout64_I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout65_I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(BitIn));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(EN));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(RST));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output34_I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output35_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output39_I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output40_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output41_I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_74 ();
 gf180mcu_fd_sc_mcu7t5v0__tieh OQPSK_PS_RCOSINE2_100 (.Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__tieh OQPSK_PS_RCOSINE2_101 (.Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__tieh OQPSK_PS_RCOSINE2_102 (.Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__tieh OQPSK_PS_RCOSINE2_103 (.Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__tieh OQPSK_PS_RCOSINE2_104 (.Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_PS_RCOSINE2_67 (.ZN(net67));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_PS_RCOSINE2_68 (.ZN(net68));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_PS_RCOSINE2_69 (.ZN(net69));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_PS_RCOSINE2_70 (.ZN(net70));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_PS_RCOSINE2_71 (.ZN(net71));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_PS_RCOSINE2_72 (.ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_PS_RCOSINE2_73 (.ZN(net73));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_PS_RCOSINE2_74 (.ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_PS_RCOSINE2_75 (.ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_PS_RCOSINE2_76 (.ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_PS_RCOSINE2_77 (.ZN(net77));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_PS_RCOSINE2_78 (.ZN(net78));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_PS_RCOSINE2_79 (.ZN(net79));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_PS_RCOSINE2_80 (.ZN(net80));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_PS_RCOSINE2_81 (.ZN(net81));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_PS_RCOSINE2_82 (.ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_PS_RCOSINE2_83 (.ZN(net83));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_PS_RCOSINE2_84 (.ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_PS_RCOSINE2_85 (.ZN(net85));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_PS_RCOSINE2_86 (.ZN(net86));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_PS_RCOSINE2_87 (.ZN(net87));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_PS_RCOSINE2_88 (.ZN(net88));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_PS_RCOSINE2_89 (.ZN(net89));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_PS_RCOSINE2_90 (.ZN(net90));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_PS_RCOSINE2_91 (.ZN(net91));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_PS_RCOSINE2_92 (.ZN(net92));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_PS_RCOSINE2_93 (.ZN(net93));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_PS_RCOSINE2_94 (.ZN(net94));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_PS_RCOSINE2_95 (.ZN(net95));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_PS_RCOSINE2_96 (.ZN(net96));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_PS_RCOSINE2_97 (.ZN(net97));
 gf180mcu_fd_sc_mcu7t5v0__tieh OQPSK_PS_RCOSINE2_98 (.Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__tieh OQPSK_PS_RCOSINE2_99 (.Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1442_ (.I(net54),
    .Z(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1443_ (.I(_1258_),
    .ZN(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1444_ (.I(_1268_),
    .Z(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1445_ (.I(net53),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1446_ (.I(_1288_),
    .Z(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1447_ (.I(_1299_),
    .Z(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1448_ (.I(net55),
    .Z(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1449_ (.I(_1321_),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1450_ (.I(_1332_),
    .Z(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1451_ (.I(net32),
    .Z(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1452_ (.I(_1354_),
    .Z(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1453_ (.I(_1365_),
    .Z(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1454_ (.A1(_1343_),
    .A2(_1376_),
    .ZN(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1455_ (.A1(_1277_),
    .A2(_1310_),
    .A3(_1387_),
    .ZN(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1456_ (.I(net34),
    .ZN(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1457_ (.A1(net35),
    .A2(_1408_),
    .ZN(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1458_ (.I(net32),
    .ZN(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1459_ (.I(_1430_),
    .Z(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1460_ (.I(net54),
    .Z(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1461_ (.I(net55),
    .Z(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1462_ (.I(net32),
    .Z(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1463_ (.A1(_0036_),
    .A2(_0047_),
    .A3(_0058_),
    .Z(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1464_ (.I0(_1441_),
    .I1(_0069_),
    .S(_1288_),
    .Z(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1465_ (.I(net53),
    .Z(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1466_ (.A1(_1258_),
    .A2(_1354_),
    .Z(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1467_ (.I(_0102_),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1468_ (.I(net34),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1469_ (.I(net35),
    .Z(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _1470_ (.A1(_0091_),
    .A2(_0113_),
    .B(_0124_),
    .C(_0135_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1471_ (.I(net54),
    .Z(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1472_ (.A1(_0157_),
    .A2(_1365_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1473_ (.I(net53),
    .Z(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1474_ (.A1(_0178_),
    .A2(net34),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1475_ (.I(net35),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1476_ (.I(_0200_),
    .Z(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1477_ (.A1(_0168_),
    .A2(_0189_),
    .B(_0211_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _1478_ (.A1(_1419_),
    .A2(_0080_),
    .B(_0146_),
    .C(_0222_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1479_ (.A1(_1397_),
    .A2(_0233_),
    .Z(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1480_ (.I(_0243_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1481_ (.I(_0254_),
    .Z(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1482_ (.I(_0265_),
    .Z(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1483_ (.I(net52),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1484_ (.I(_0286_),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1485_ (.I(_0297_),
    .Z(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1486_ (.I(net51),
    .Z(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1487_ (.I(_0318_),
    .Z(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1488_ (.I(net50),
    .Z(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1489_ (.I(_0340_),
    .Z(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1490_ (.I(net38),
    .Z(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1491_ (.I(_0361_),
    .Z(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1492_ (.I(_0371_),
    .Z(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _1493_ (.A1(_0329_),
    .A2(_0351_),
    .A3(_0382_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1494_ (.A1(_0308_),
    .A2(_0393_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1495_ (.I(net38),
    .Z(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1496_ (.A1(_0340_),
    .A2(_0414_),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1497_ (.I(net50),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1498_ (.I(_0436_),
    .Z(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1499_ (.I(_0447_),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1500_ (.I(_0318_),
    .Z(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1501_ (.I(_0286_),
    .Z(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1502_ (.I(_0361_),
    .Z(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _1503_ (.A1(_0468_),
    .A2(_0479_),
    .A3(_0489_),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1504_ (.A1(_0457_),
    .A2(_0500_),
    .ZN(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1505_ (.I(net49),
    .Z(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1506_ (.I(net40),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1507_ (.I(_0532_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1508_ (.A1(_0521_),
    .A2(_0542_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1509_ (.A1(_0425_),
    .A2(_0511_),
    .B(_0553_),
    .ZN(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1510_ (.I(net49),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1511_ (.I(_0532_),
    .Z(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _1512_ (.A1(_0569_),
    .A2(_0577_),
    .A3(_0393_),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1513_ (.I(net40),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1514_ (.I(_0592_),
    .Z(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1515_ (.I(_0436_),
    .Z(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1516_ (.I(_0361_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1517_ (.A1(_0468_),
    .A2(_0600_),
    .ZN(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1518_ (.A1(_0599_),
    .A2(_0601_),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1519_ (.I(net49),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1520_ (.A1(_0598_),
    .A2(_0602_),
    .B(_0603_),
    .ZN(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1521_ (.A1(_0404_),
    .A2(_0562_),
    .A3(_0585_),
    .A4(_0604_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1522_ (.I(_0605_),
    .Z(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1523_ (.I(\p_shaping_I.bit_in_1 ),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1524_ (.I(_0606_),
    .Z(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1525_ (.I(_0607_),
    .Z(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1526_ (.I(_0243_),
    .Z(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1527_ (.I(\p_shaping_I.bit_in ),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1528_ (.I(_0610_),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1529_ (.I(net63),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1530_ (.A1(\p_shaping_I.ctl_1 ),
    .A2(_0612_),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1531_ (.A1(_0611_),
    .A2(_0612_),
    .B(_0613_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1532_ (.A1(_0609_),
    .A2(_0614_),
    .ZN(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1533_ (.A1(_0608_),
    .A2(_0609_),
    .B(_0615_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1534_ (.I(\p_shaping_Q.bit_in_1 ),
    .Z(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1535_ (.I(_0616_),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1536_ (.I(_0617_),
    .Z(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1537_ (.I(\Reg_Delay_Q.Out ),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1538_ (.A1(net62),
    .A2(\p_shaping_Q.ctl_1 ),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1539_ (.A1(_0612_),
    .A2(_0619_),
    .B(_0620_),
    .ZN(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1540_ (.A1(net47),
    .A2(_0621_),
    .ZN(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1541_ (.A1(_0618_),
    .A2(net47),
    .B(_0622_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1542_ (.I(_0612_),
    .ZN(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1543_ (.A1(_0623_),
    .A2(net42),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1544_ (.A1(_0623_),
    .A2(net47),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1545_ (.I(_0585_),
    .Z(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1546_ (.I(_0286_),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1547_ (.I(_0625_),
    .Z(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1548_ (.I(net38),
    .ZN(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1549_ (.I(_0627_),
    .Z(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1550_ (.I(_0628_),
    .Z(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1551_ (.A1(_0626_),
    .A2(_0629_),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1552_ (.I(_0630_),
    .Z(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1553_ (.I(net51),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1554_ (.I(_0632_),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1555_ (.I(_0633_),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1556_ (.I(_0414_),
    .Z(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _1557_ (.A1(_0634_),
    .A2(_0479_),
    .A3(_0635_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1558_ (.I(_0457_),
    .Z(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1559_ (.A1(_0631_),
    .A2(_0636_),
    .B(_0637_),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1560_ (.I(_0577_),
    .Z(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1561_ (.I(_0286_),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1562_ (.I(_0640_),
    .Z(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1563_ (.I(_0371_),
    .Z(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1564_ (.I(net50),
    .Z(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1565_ (.I(_0643_),
    .Z(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1566_ (.A1(_0641_),
    .A2(_0642_),
    .B(_0644_),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1567_ (.I(_0645_),
    .Z(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1568_ (.I(_0633_),
    .Z(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1569_ (.I(_0371_),
    .Z(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1570_ (.I(_0648_),
    .Z(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1571_ (.A1(_0647_),
    .A2(_0649_),
    .B(_0645_),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1572_ (.I(_0632_),
    .Z(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1573_ (.A1(_0651_),
    .A2(_0640_),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1574_ (.I(_0652_),
    .Z(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1575_ (.A1(_0639_),
    .A2(_0646_),
    .B1(_0650_),
    .B2(_0653_),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1576_ (.I(_0521_),
    .Z(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1577_ (.I(_0655_),
    .Z(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1578_ (.A1(_0638_),
    .A2(_0654_),
    .B(_0656_),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1579_ (.A1(_0468_),
    .A2(_0629_),
    .B(_0599_),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1580_ (.I(_0489_),
    .Z(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1581_ (.I(_0659_),
    .Z(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1582_ (.A1(net51),
    .A2(net52),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1583_ (.I(_0661_),
    .Z(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1584_ (.I(_0662_),
    .Z(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1585_ (.I(_0643_),
    .Z(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1586_ (.I(_0664_),
    .Z(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _1587_ (.A1(_0660_),
    .A2(_0663_),
    .B(_0500_),
    .C(_0665_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1588_ (.A1(_0658_),
    .A2(_0666_),
    .B(_0553_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1589_ (.A1(_0624_),
    .A2(_0657_),
    .A3(_0667_),
    .Z(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1590_ (.A1(\p_shaping_Q.counter[1] ),
    .A2(\p_shaping_Q.counter[0] ),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1591_ (.I(_0669_),
    .ZN(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1592_ (.I(_0670_),
    .Z(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1593_ (.I(_0671_),
    .Z(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1594_ (.I(net40),
    .Z(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1595_ (.I(_0673_),
    .Z(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1596_ (.I(net52),
    .Z(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1597_ (.A1(_0651_),
    .A2(_0675_),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1598_ (.I(_0632_),
    .Z(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1599_ (.I(_0361_),
    .Z(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1600_ (.A1(_0677_),
    .A2(_0678_),
    .Z(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1601_ (.A1(_0351_),
    .A2(_0676_),
    .A3(_0679_),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1602_ (.I(_0675_),
    .Z(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1603_ (.I(_0340_),
    .Z(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _1604_ (.A1(_0681_),
    .A2(_0682_),
    .A3(_0635_),
    .Z(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _1605_ (.A1(_0318_),
    .A2(_0675_),
    .A3(_0340_),
    .A4(_0414_),
    .Z(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _1606_ (.A1(net49),
    .A2(_0684_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _1607_ (.A1(_0521_),
    .A2(_0680_),
    .A3(_0683_),
    .B(_0685_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1608_ (.I(_0600_),
    .Z(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1609_ (.A1(_0634_),
    .A2(_0681_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1610_ (.A1(_0635_),
    .A2(_0652_),
    .B(_0682_),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1611_ (.A1(_0687_),
    .A2(_0688_),
    .B(_0689_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1612_ (.I(net50),
    .Z(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1613_ (.I(_0632_),
    .Z(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1614_ (.A1(_0692_),
    .A2(_0371_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1615_ (.A1(_0691_),
    .A2(_0661_),
    .A3(_0693_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1616_ (.A1(_0521_),
    .A2(_0592_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1617_ (.A1(_0694_),
    .A2(_0695_),
    .Z(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1618_ (.A1(_0318_),
    .A2(_0628_),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1619_ (.I0(_0457_),
    .I1(_0658_),
    .S(_0697_),
    .Z(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1620_ (.I(_0685_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _1621_ (.A1(_0674_),
    .A2(_0686_),
    .B1(_0690_),
    .B2(_0696_),
    .C1(_0698_),
    .C2(_0699_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1622_ (.I(\p_shaping_Q.counter[1] ),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1623_ (.I(_0701_),
    .Z(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1624_ (.I(_0664_),
    .Z(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1625_ (.I(_0676_),
    .Z(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _1626_ (.A1(_0703_),
    .A2(_0674_),
    .A3(_0704_),
    .B(_0655_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1627_ (.I(_0542_),
    .Z(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1628_ (.I(_0682_),
    .Z(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1629_ (.I(_0633_),
    .Z(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1630_ (.I(_0628_),
    .Z(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1631_ (.A1(_0708_),
    .A2(_0709_),
    .B(_0641_),
    .ZN(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1632_ (.A1(_0651_),
    .A2(_0675_),
    .B(_0414_),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1633_ (.A1(_0664_),
    .A2(_0711_),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1634_ (.A1(_0651_),
    .A2(_0640_),
    .Z(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1635_ (.I(_0713_),
    .Z(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1636_ (.A1(_0707_),
    .A2(_0710_),
    .B1(_0712_),
    .B2(_0714_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1637_ (.A1(net37),
    .A2(net36),
    .Z(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1638_ (.A1(_0692_),
    .A2(_0678_),
    .B(_0643_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1639_ (.A1(_0382_),
    .A2(_0716_),
    .B(_0717_),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1640_ (.I(_0532_),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1641_ (.I(_0447_),
    .Z(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1642_ (.A1(_0687_),
    .A2(_0704_),
    .B(_0720_),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1643_ (.A1(_0719_),
    .A2(_0721_),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1644_ (.I(_0569_),
    .Z(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _1645_ (.A1(_0706_),
    .A2(_0715_),
    .B1(_0718_),
    .B2(_0722_),
    .C(_0723_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1646_ (.A1(_0705_),
    .A2(_0724_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1647_ (.A1(_0702_),
    .A2(_0725_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1648_ (.A1(_0700_),
    .A2(_0726_),
    .Z(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1649_ (.A1(_0672_),
    .A2(_0727_),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1650_ (.A1(_0668_),
    .A2(_0728_),
    .Z(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1651_ (.I(_0729_),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1652_ (.I(_0702_),
    .Z(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1653_ (.I(_0730_),
    .Z(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1654_ (.I(_0706_),
    .Z(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1655_ (.I(_0603_),
    .Z(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _1656_ (.I(_0684_),
    .Z(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1657_ (.I(_0457_),
    .Z(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1658_ (.A1(_0735_),
    .A2(_0714_),
    .A3(_0693_),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1659_ (.A1(_0655_),
    .A2(_0683_),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1660_ (.A1(_0733_),
    .A2(_0734_),
    .B1(_0736_),
    .B2(_0737_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1661_ (.I(_0329_),
    .Z(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1662_ (.I(_0626_),
    .Z(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1663_ (.A1(_0739_),
    .A2(_0740_),
    .B(_0659_),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1664_ (.I(_0691_),
    .Z(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1665_ (.I(_0742_),
    .Z(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _1666_ (.A1(_0660_),
    .A2(_0653_),
    .B(_0741_),
    .C(_0743_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1667_ (.A1(_0694_),
    .A2(_0695_),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1668_ (.I(_0682_),
    .Z(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1669_ (.A1(_0647_),
    .A2(_0659_),
    .B(_0746_),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1670_ (.I(_0697_),
    .Z(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1671_ (.I0(_0703_),
    .I1(_0747_),
    .S(_0748_),
    .Z(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_4 _1672_ (.A1(_0732_),
    .A2(_0738_),
    .B1(_0744_),
    .B2(_0745_),
    .C1(_0749_),
    .C2(_0685_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _1673_ (.A1(_0731_),
    .A2(_0750_),
    .A3(_0725_),
    .B1(_0728_),
    .B2(_0668_),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1674_ (.I(\Reg_Delay_Q.Out ),
    .Z(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1675_ (.A1(_0752_),
    .A2(_0668_),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1676_ (.I(_0553_),
    .Z(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1677_ (.I(_0711_),
    .Z(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1678_ (.A1(_0709_),
    .A2(_0662_),
    .B(_0599_),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1679_ (.A1(_0755_),
    .A2(_0756_),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1680_ (.I(_0723_),
    .Z(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1681_ (.I(_0627_),
    .Z(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1682_ (.I(_0759_),
    .Z(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1683_ (.A1(_0647_),
    .A2(_0760_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1684_ (.A1(_0677_),
    .A2(_0297_),
    .A3(_0600_),
    .Z(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1685_ (.I(_0762_),
    .Z(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1686_ (.I(_0640_),
    .Z(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1687_ (.A1(_0764_),
    .A2(_0642_),
    .B(_0708_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1688_ (.I0(_0761_),
    .I1(_0763_),
    .I2(_0765_),
    .I3(_0688_),
    .S0(_0719_),
    .S1(_0735_),
    .Z(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1689_ (.A1(_0758_),
    .A2(_0766_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _1690_ (.A1(_0754_),
    .A2(_0650_),
    .A3(_0757_),
    .B(_0767_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1691_ (.A1(_0753_),
    .A2(_0768_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1692_ (.I(_0569_),
    .Z(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1693_ (.I(_0770_),
    .Z(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1694_ (.A1(_0329_),
    .A2(_0709_),
    .B(_0626_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _1695_ (.A1(_0720_),
    .A2(_0772_),
    .B(_0636_),
    .C(_0630_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1696_ (.A1(_0425_),
    .A2(_0652_),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1697_ (.A1(_0673_),
    .A2(_0774_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _1698_ (.A1(_0703_),
    .A2(_0748_),
    .B1(_0773_),
    .B2(_0674_),
    .C(_0775_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _1699_ (.A1(_0692_),
    .A2(_0643_),
    .A3(_0678_),
    .Z(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1700_ (.I(_0628_),
    .Z(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1701_ (.A1(_0778_),
    .A2(_0676_),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _1702_ (.A1(_0329_),
    .A2(_0626_),
    .A3(_0629_),
    .B(_0542_),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1703_ (.I(_0716_),
    .Z(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1704_ (.A1(_0648_),
    .A2(_0781_),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _1705_ (.A1(_0742_),
    .A2(_0779_),
    .B(_0780_),
    .C(_0782_),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _1706_ (.A1(_0674_),
    .A2(_0777_),
    .B(_0783_),
    .C(_0723_),
    .ZN(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1707_ (.A1(_0771_),
    .A2(_0776_),
    .B(_0784_),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1708_ (.A1(_0616_),
    .A2(_0750_),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1709_ (.A1(_0785_),
    .A2(_0786_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1710_ (.I(\p_shaping_Q.counter[1] ),
    .Z(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1711_ (.I(\p_shaping_Q.bit_in_2 ),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1712_ (.I(_0692_),
    .Z(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _1713_ (.A1(_0297_),
    .A2(_0600_),
    .Z(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _1714_ (.A1(_0790_),
    .A2(_0778_),
    .B(_0791_),
    .C(_0644_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1715_ (.I(_0592_),
    .Z(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1716_ (.A1(_0792_),
    .A2(_0756_),
    .B(_0793_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1717_ (.I(_0447_),
    .Z(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1718_ (.A1(_0795_),
    .A2(_0577_),
    .A3(_0662_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _1719_ (.A1(_0708_),
    .A2(_0641_),
    .B(_0644_),
    .C(_0648_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1720_ (.A1(_0425_),
    .A2(_0713_),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1721_ (.A1(_0797_),
    .A2(_0798_),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1722_ (.A1(_0598_),
    .A2(_0684_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1723_ (.A1(_0603_),
    .A2(_0800_),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _1724_ (.A1(_0655_),
    .A2(_0794_),
    .A3(_0796_),
    .B1(_0799_),
    .B2(_0801_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1725_ (.A1(_0789_),
    .A2(_0705_),
    .A3(_0724_),
    .A4(_0802_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1726_ (.I(\p_shaping_Q.bit_in_2 ),
    .Z(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1727_ (.I(_0705_),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1728_ (.I(_0673_),
    .Z(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1729_ (.I(_0806_),
    .Z(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1730_ (.I(_0807_),
    .Z(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1731_ (.I(_0735_),
    .Z(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1732_ (.I(_0625_),
    .Z(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1733_ (.A1(_0790_),
    .A2(_0642_),
    .B(_0810_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1734_ (.I(_0707_),
    .Z(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1735_ (.I(_0676_),
    .Z(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1736_ (.A1(_0812_),
    .A2(_0813_),
    .A3(_0755_),
    .Z(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1737_ (.A1(_0809_),
    .A2(_0811_),
    .B(_0814_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1738_ (.I(_0599_),
    .Z(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1739_ (.I(_0816_),
    .Z(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1740_ (.I(_0629_),
    .Z(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1741_ (.A1(_0818_),
    .A2(_0714_),
    .ZN(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1742_ (.I(_0806_),
    .Z(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1743_ (.A1(_0817_),
    .A2(_0819_),
    .B(_0718_),
    .C(_0820_),
    .ZN(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1744_ (.I(_0656_),
    .Z(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1745_ (.A1(_0808_),
    .A2(_0815_),
    .B(_0821_),
    .C(_0822_),
    .ZN(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1746_ (.A1(_0797_),
    .A2(_0798_),
    .Z(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1747_ (.A1(_0793_),
    .A2(_0734_),
    .B(_0723_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1748_ (.A1(_0382_),
    .A2(_0781_),
    .B(_0351_),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1749_ (.A1(_0650_),
    .A2(_0826_),
    .B(_0732_),
    .ZN(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1750_ (.I(_0733_),
    .Z(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1751_ (.A1(_0828_),
    .A2(_0796_),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1752_ (.A1(_0824_),
    .A2(_0825_),
    .B1(_0827_),
    .B2(_0829_),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1753_ (.A1(_0804_),
    .A2(_0805_),
    .A3(_0823_),
    .B(_0830_),
    .ZN(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1754_ (.A1(_0788_),
    .A2(_0803_),
    .A3(_0831_),
    .Z(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1755_ (.A1(_0787_),
    .A2(_0832_),
    .Z(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1756_ (.A1(_0787_),
    .A2(_0832_),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1757_ (.A1(_0670_),
    .A2(_0833_),
    .A3(_0834_),
    .ZN(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1758_ (.A1(_0769_),
    .A2(_0835_),
    .Z(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1759_ (.A1(_0751_),
    .A2(_0836_),
    .Z(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1760_ (.A1(_0769_),
    .A2(_0835_),
    .B(_0834_),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _1761_ (.A1(_0585_),
    .A2(_0657_),
    .A3(_0667_),
    .ZN(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1762_ (.A1(_0839_),
    .A2(_0768_),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1763_ (.A1(_0752_),
    .A2(_0840_),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1764_ (.I(_0793_),
    .Z(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1765_ (.A1(_0743_),
    .A2(_0710_),
    .B(_0842_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1766_ (.I(_0308_),
    .Z(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1767_ (.A1(_0844_),
    .A2(_0817_),
    .A3(_0748_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1768_ (.A1(_0656_),
    .A2(_0843_),
    .A3(_0845_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1769_ (.A1(_0649_),
    .A2(_0652_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _1770_ (.A1(_0677_),
    .A2(_0625_),
    .A3(_0759_),
    .B(_0447_),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1771_ (.I(_0848_),
    .Z(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1772_ (.A1(_0637_),
    .A2(_0763_),
    .B1(_0847_),
    .B2(_0849_),
    .C(_0639_),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1773_ (.I(_0592_),
    .Z(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1774_ (.I(_0851_),
    .Z(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1775_ (.A1(_0760_),
    .A2(_0662_),
    .ZN(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1776_ (.I(_0760_),
    .Z(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1777_ (.A1(_0790_),
    .A2(_0764_),
    .Z(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1778_ (.A1(_0854_),
    .A2(_0855_),
    .B(_0665_),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1779_ (.A1(_0852_),
    .A2(_0853_),
    .A3(_0856_),
    .ZN(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1780_ (.A1(_0850_),
    .A2(_0857_),
    .Z(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1781_ (.A1(_0822_),
    .A2(_0858_),
    .Z(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1782_ (.A1(_0846_),
    .A2(_0859_),
    .Z(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1783_ (.A1(_0841_),
    .A2(_0860_),
    .Z(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1784_ (.I(_0669_),
    .Z(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1785_ (.I(\p_shaping_Q.bit_in_1 ),
    .Z(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _1786_ (.A1(_0758_),
    .A2(_0776_),
    .B(_0784_),
    .C(_0700_),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1787_ (.A1(_0863_),
    .A2(_0864_),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1788_ (.A1(_0625_),
    .A2(_0759_),
    .B(_0677_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1789_ (.A1(_0634_),
    .A2(_0382_),
    .B(_0681_),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _1790_ (.A1(_0795_),
    .A2(_0866_),
    .B1(_0867_),
    .B2(_0848_),
    .C(_0577_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1791_ (.I(_0634_),
    .Z(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1792_ (.A1(_0869_),
    .A2(_0764_),
    .A3(_0664_),
    .A4(_0778_),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1793_ (.A1(_0308_),
    .A2(_0720_),
    .A3(_0679_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1794_ (.A1(_0870_),
    .A2(_0871_),
    .B(_0851_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _1795_ (.A1(_0770_),
    .A2(_0868_),
    .A3(_0872_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1796_ (.A1(_0810_),
    .A2(_0777_),
    .B(_0673_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1797_ (.A1(_0603_),
    .A2(_0874_),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1798_ (.A1(_0746_),
    .A2(_0765_),
    .B(_0826_),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1799_ (.A1(_0875_),
    .A2(_0876_),
    .Z(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1800_ (.A1(_0873_),
    .A2(_0877_),
    .Z(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1801_ (.A1(_0619_),
    .A2(_0620_),
    .Z(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1802_ (.A1(_0605_),
    .A2(_0879_),
    .Z(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1803_ (.A1(_0878_),
    .A2(_0880_),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1804_ (.A1(_0865_),
    .A2(_0881_),
    .Z(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1805_ (.A1(_0705_),
    .A2(_0724_),
    .B(_0802_),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1806_ (.I(_0883_),
    .Z(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1807_ (.A1(_0804_),
    .A2(_0884_),
    .Z(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1808_ (.A1(_0569_),
    .A2(_0598_),
    .ZN(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1809_ (.I(_0886_),
    .Z(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1810_ (.I0(_0631_),
    .I1(_0741_),
    .S(_0816_),
    .Z(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1811_ (.I(_0425_),
    .Z(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1812_ (.A1(_0869_),
    .A2(_0764_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1813_ (.A1(_0889_),
    .A2(_0890_),
    .ZN(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1814_ (.A1(_0479_),
    .A2(_0489_),
    .B(_0691_),
    .ZN(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1815_ (.A1(_0708_),
    .A2(_0641_),
    .B(_0648_),
    .ZN(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1816_ (.A1(_0793_),
    .A2(_0893_),
    .Z(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1817_ (.A1(_0762_),
    .A2(_0711_),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1818_ (.A1(_0740_),
    .A2(_0707_),
    .A3(_0697_),
    .B1(_0797_),
    .B2(_0895_),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _1819_ (.A1(_0891_),
    .A2(_0892_),
    .A3(_0894_),
    .B1(_0896_),
    .B2(_0639_),
    .ZN(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _1820_ (.A1(_0887_),
    .A2(_0888_),
    .B1(_0897_),
    .B2(_0758_),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1821_ (.I(_0898_),
    .Z(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1822_ (.A1(_0804_),
    .A2(_0884_),
    .A3(_0899_),
    .B(_0788_),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1823_ (.A1(_0885_),
    .A2(_0899_),
    .B(_0900_),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1824_ (.A1(_0882_),
    .A2(_0901_),
    .ZN(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1825_ (.A1(_0862_),
    .A2(_0902_),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _1826_ (.A1(_0838_),
    .A2(_0861_),
    .A3(_0903_),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1827_ (.A1(_0837_),
    .A2(_0904_),
    .Z(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1828_ (.I(_0905_),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1829_ (.A1(_0882_),
    .A2(_0901_),
    .ZN(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _1830_ (.A1(_0862_),
    .A2(_0861_),
    .A3(_0902_),
    .B(_0906_),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1831_ (.A1(_0840_),
    .A2(_0860_),
    .B(_0752_),
    .ZN(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1832_ (.I(_0733_),
    .Z(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1833_ (.A1(_0633_),
    .A2(_0297_),
    .B(_0678_),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1834_ (.I(_0910_),
    .Z(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1835_ (.A1(_0817_),
    .A2(_0911_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1836_ (.A1(_0740_),
    .A2(_0649_),
    .B(_0637_),
    .ZN(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1837_ (.A1(_0742_),
    .A2(_0659_),
    .Z(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1838_ (.A1(_0914_),
    .A2(_0813_),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1839_ (.A1(_0818_),
    .A2(_0704_),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1840_ (.A1(_0813_),
    .A2(_0913_),
    .B(_0915_),
    .C(_0916_),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1841_ (.A1(_0843_),
    .A2(_0912_),
    .B1(_0917_),
    .B2(_0852_),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1842_ (.A1(_0665_),
    .A2(_0649_),
    .A3(_0781_),
    .ZN(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1843_ (.A1(_0646_),
    .A2(_0663_),
    .B(_0706_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1844_ (.A1(_0919_),
    .A2(_0920_),
    .B(_0404_),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1845_ (.A1(_0656_),
    .A2(_0921_),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1846_ (.A1(_0909_),
    .A2(_0918_),
    .B(_0922_),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1847_ (.A1(_0908_),
    .A2(_0923_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1848_ (.I(_0788_),
    .Z(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1849_ (.A1(_0351_),
    .A2(_0866_),
    .ZN(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1850_ (.A1(_0479_),
    .A2(_0759_),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1851_ (.A1(_0635_),
    .A2(_0716_),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1852_ (.A1(_0927_),
    .A2(_0928_),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1853_ (.A1(_0926_),
    .A2(_0929_),
    .Z(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1854_ (.A1(_0748_),
    .A2(_0911_),
    .B(_0746_),
    .C(_0704_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1855_ (.A1(_0869_),
    .A2(_0687_),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1856_ (.A1(_0790_),
    .A2(_0810_),
    .B(_0778_),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1857_ (.A1(_0795_),
    .A2(_0932_),
    .A3(_0933_),
    .B(_0851_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1858_ (.A1(_0468_),
    .A2(_0489_),
    .B(_0691_),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1859_ (.A1(_0810_),
    .A2(_0642_),
    .B(_0935_),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1860_ (.A1(_0792_),
    .A2(_0895_),
    .B(_0936_),
    .C(_0719_),
    .ZN(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1861_ (.A1(_0931_),
    .A2(_0934_),
    .B(_0937_),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _1862_ (.A1(_0886_),
    .A2(_0930_),
    .B1(_0938_),
    .B2(_0770_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1863_ (.A1(_0884_),
    .A2(_0899_),
    .B(\p_shaping_Q.bit_in_2 ),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1864_ (.A1(_0939_),
    .A2(_0940_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1865_ (.A1(_0605_),
    .A2(_0879_),
    .ZN(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1866_ (.A1(_0687_),
    .A2(_0713_),
    .ZN(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1867_ (.A1(_0853_),
    .A2(_0943_),
    .B(_0816_),
    .ZN(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1868_ (.A1(_0747_),
    .A2(_0944_),
    .B(_0825_),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1869_ (.A1(_0697_),
    .A2(_0910_),
    .B(_0746_),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1870_ (.A1(_0598_),
    .A2(_0718_),
    .Z(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1871_ (.A1(_0542_),
    .A2(_0892_),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1872_ (.A1(_0795_),
    .A2(_0811_),
    .B(_0948_),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _1873_ (.A1(_0946_),
    .A2(_0947_),
    .B(_0949_),
    .C(_0770_),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1874_ (.A1(_0942_),
    .A2(_0945_),
    .A3(_0950_),
    .Z(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1875_ (.A1(_0864_),
    .A2(_0878_),
    .B(_0616_),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1876_ (.A1(_0951_),
    .A2(_0952_),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1877_ (.A1(_0925_),
    .A2(_0941_),
    .B(_0953_),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1878_ (.A1(_0788_),
    .A2(_0941_),
    .A3(_0953_),
    .Z(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _1879_ (.A1(_0669_),
    .A2(_0924_),
    .A3(_0954_),
    .A4(_0955_),
    .Z(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _1880_ (.A1(_0862_),
    .A2(_0954_),
    .A3(_0955_),
    .B(_0924_),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1881_ (.A1(_0956_),
    .A2(_0957_),
    .ZN(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1882_ (.A1(_0862_),
    .A2(_0861_),
    .A3(_0902_),
    .Z(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1883_ (.I(_0669_),
    .Z(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1884_ (.A1(_0960_),
    .A2(_0902_),
    .B(_0861_),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1885_ (.A1(_0838_),
    .A2(_0959_),
    .A3(_0961_),
    .Z(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1886_ (.A1(_0837_),
    .A2(_0904_),
    .B(_0962_),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1887_ (.A1(_0907_),
    .A2(_0958_),
    .A3(_0963_),
    .Z(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1888_ (.I(_0964_),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1889_ (.I(_0955_),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1890_ (.A1(_0965_),
    .A2(_0956_),
    .ZN(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1891_ (.I(_0743_),
    .Z(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1892_ (.A1(_0818_),
    .A2(_0653_),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1893_ (.I(_0943_),
    .Z(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1894_ (.A1(_0968_),
    .A2(_0969_),
    .ZN(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1895_ (.I(_0665_),
    .Z(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1896_ (.A1(_0971_),
    .A2(_0855_),
    .ZN(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1897_ (.A1(_0967_),
    .A2(_0970_),
    .B1(_0972_),
    .B2(_0791_),
    .C(_0754_),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1898_ (.I(_0732_),
    .Z(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1899_ (.I(_0693_),
    .Z(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1900_ (.A1(_0637_),
    .A2(_0975_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1901_ (.A1(_0739_),
    .A2(_0976_),
    .ZN(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1902_ (.A1(_0971_),
    .A2(_0975_),
    .A3(_0819_),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1903_ (.A1(_0974_),
    .A2(_0977_),
    .B1(_0978_),
    .B2(_0948_),
    .C(_0828_),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1904_ (.A1(_0973_),
    .A2(_0979_),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1905_ (.A1(_0828_),
    .A2(_0858_),
    .B(_0846_),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1906_ (.A1(_0839_),
    .A2(_0768_),
    .A3(_0981_),
    .A4(_0923_),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1907_ (.A1(_0752_),
    .A2(_0982_),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1908_ (.A1(_0980_),
    .A2(_0983_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1909_ (.I(_0789_),
    .Z(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1910_ (.A1(_0884_),
    .A2(_0899_),
    .A3(_0939_),
    .ZN(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1911_ (.A1(_0694_),
    .A2(_0756_),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1912_ (.A1(_0816_),
    .A2(_0855_),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1913_ (.A1(_0681_),
    .A2(_0709_),
    .B(_0644_),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1914_ (.A1(_0308_),
    .A2(_0760_),
    .B(_0869_),
    .ZN(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _1915_ (.A1(_0867_),
    .A2(_0849_),
    .B1(_0989_),
    .B2(_0990_),
    .C(_0851_),
    .ZN(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _1916_ (.A1(_0806_),
    .A2(_0935_),
    .A3(_0988_),
    .B(_0991_),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _1917_ (.A1(_0887_),
    .A2(_0987_),
    .B1(_0992_),
    .B2(_0758_),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1918_ (.I(_0993_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1919_ (.A1(_0985_),
    .A2(_0986_),
    .A3(_0994_),
    .Z(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1920_ (.A1(_0985_),
    .A2(_0986_),
    .B(_0994_),
    .ZN(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1921_ (.A1(_0873_),
    .A2(_0877_),
    .A3(_0945_),
    .A4(_0950_),
    .Z(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1922_ (.A1(_0864_),
    .A2(_0997_),
    .B(_0616_),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1923_ (.A1(_0854_),
    .A2(_0890_),
    .B(_0772_),
    .C(_0812_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1924_ (.A1(_0761_),
    .A2(_0943_),
    .B(_0842_),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _1925_ (.A1(_0807_),
    .A2(_0734_),
    .B1(_0999_),
    .B2(_1000_),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1926_ (.A1(_0717_),
    .A2(_0679_),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1927_ (.A1(_0739_),
    .A2(_0703_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1928_ (.A1(_0735_),
    .A2(_0636_),
    .Z(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1929_ (.A1(_0806_),
    .A2(_0890_),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1930_ (.A1(_0842_),
    .A2(_1002_),
    .A3(_1003_),
    .B1(_1004_),
    .B2(_1005_),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1931_ (.A1(_0771_),
    .A2(_1006_),
    .Z(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1932_ (.A1(_0828_),
    .A2(_1001_),
    .B(_1007_),
    .C(_0880_),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1933_ (.A1(_0998_),
    .A2(_1008_),
    .Z(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1934_ (.A1(_0701_),
    .A2(_0995_),
    .A3(_0996_),
    .B(_1009_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1935_ (.A1(_0701_),
    .A2(_1009_),
    .A3(_0995_),
    .A4(_0996_),
    .Z(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1936_ (.A1(_0671_),
    .A2(_1010_),
    .A3(_1011_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1937_ (.A1(_0984_),
    .A2(_1012_),
    .ZN(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _1938_ (.A1(_0966_),
    .A2(_1013_),
    .ZN(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1939_ (.A1(_0956_),
    .A2(_0957_),
    .B(_0907_),
    .ZN(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1940_ (.A1(_0907_),
    .A2(_0956_),
    .A3(_0957_),
    .Z(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _1941_ (.A1(_0837_),
    .A2(_0904_),
    .B(_1016_),
    .C(_0962_),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1942_ (.A1(_1015_),
    .A2(_1017_),
    .Z(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1943_ (.A1(_1014_),
    .A2(_1018_),
    .Z(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1944_ (.I(_1019_),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1945_ (.A1(_0730_),
    .A2(_1009_),
    .A3(_0995_),
    .A4(_0996_),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1946_ (.A1(_0672_),
    .A2(_0984_),
    .A3(_1010_),
    .A4(_1011_),
    .Z(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1947_ (.A1(_1020_),
    .A2(_1021_),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1948_ (.I(_0853_),
    .Z(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1949_ (.A1(_1023_),
    .A2(_0892_),
    .B(_0820_),
    .C(_0914_),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1950_ (.I(_0852_),
    .Z(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1951_ (.A1(_0817_),
    .A2(_0631_),
    .A3(_0636_),
    .B(_0976_),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1952_ (.A1(_0971_),
    .A2(_0854_),
    .B(_0852_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1953_ (.A1(_1025_),
    .A2(_1026_),
    .B(_1027_),
    .ZN(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1954_ (.I(_0909_),
    .Z(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1955_ (.A1(_0685_),
    .A2(_1024_),
    .B1(_1028_),
    .B2(_1029_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1956_ (.I(\Reg_Delay_Q.Out ),
    .Z(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1957_ (.A1(_0980_),
    .A2(_0982_),
    .B(_1031_),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1958_ (.A1(_1030_),
    .A2(_1032_),
    .Z(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _1959_ (.A1(_0883_),
    .A2(_0898_),
    .A3(_0939_),
    .A4(_0993_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1960_ (.A1(_0601_),
    .A2(_0736_),
    .B(_0694_),
    .ZN(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1961_ (.A1(_0690_),
    .A2(_0989_),
    .B(_0842_),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1962_ (.A1(_0807_),
    .A2(_1035_),
    .B(_1036_),
    .ZN(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1963_ (.A1(_0707_),
    .A2(_0763_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1964_ (.A1(_0812_),
    .A2(_0968_),
    .B(_1038_),
    .ZN(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1965_ (.A1(_0887_),
    .A2(_1039_),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1966_ (.A1(_0909_),
    .A2(_1037_),
    .B(_1040_),
    .ZN(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1967_ (.A1(_0985_),
    .A2(_1034_),
    .A3(_1041_),
    .Z(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1968_ (.A1(_0985_),
    .A2(_1034_),
    .B(_1041_),
    .ZN(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1969_ (.I(_0880_),
    .Z(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1970_ (.A1(_0873_),
    .A2(_0877_),
    .A3(_0945_),
    .A4(_0950_),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1971_ (.I(_0646_),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1972_ (.A1(_0819_),
    .A2(_0911_),
    .B(_0743_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1973_ (.A1(_1046_),
    .A2(_1047_),
    .B(_0639_),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1974_ (.A1(_0688_),
    .A2(_0849_),
    .B(_0989_),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1975_ (.A1(_0740_),
    .A2(_0742_),
    .A3(_0693_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _1976_ (.A1(_0720_),
    .A2(_0755_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1977_ (.A1(_1050_),
    .A2(_1051_),
    .B(_0706_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1978_ (.A1(_0719_),
    .A2(_1050_),
    .A3(_1051_),
    .Z(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1979_ (.A1(_1049_),
    .A2(_1052_),
    .B(_0733_),
    .C(_1053_),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1980_ (.A1(_0909_),
    .A2(_1048_),
    .B(_1054_),
    .C(\p_shaping_Q.bit_in_1 ),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1981_ (.A1(_0617_),
    .A2(_1045_),
    .B(_1055_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1982_ (.I(_1056_),
    .Z(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1983_ (.A1(_1049_),
    .A2(_1052_),
    .B(_1053_),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1984_ (.I0(_1058_),
    .I1(_1048_),
    .S(_0822_),
    .Z(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1985_ (.A1(_0863_),
    .A2(_0997_),
    .B(_1059_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1986_ (.A1(_1044_),
    .A2(_1055_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1987_ (.A1(_1044_),
    .A2(_1057_),
    .B1(_1060_),
    .B2(_1061_),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1988_ (.A1(_0702_),
    .A2(_1042_),
    .A3(_1043_),
    .A4(_1062_),
    .Z(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1989_ (.A1(_0702_),
    .A2(_1042_),
    .A3(_1043_),
    .B(_1062_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1990_ (.A1(_0671_),
    .A2(_1063_),
    .A3(_1064_),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1991_ (.A1(_1033_),
    .A2(_1065_),
    .Z(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1992_ (.A1(_1022_),
    .A2(_1066_),
    .Z(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1993_ (.A1(_0966_),
    .A2(_1013_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1994_ (.A1(_1014_),
    .A2(_1018_),
    .B(_1068_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1995_ (.A1(_1067_),
    .A2(_1069_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1996_ (.I(_1070_),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1997_ (.A1(_1033_),
    .A2(_1065_),
    .B(_1063_),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1998_ (.A1(_0980_),
    .A2(_0982_),
    .A3(_1030_),
    .Z(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _1999_ (.A1(_1031_),
    .A2(_1072_),
    .Z(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2000_ (.I(_1025_),
    .Z(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2001_ (.I(_0818_),
    .Z(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2002_ (.A1(_1075_),
    .A2(_0781_),
    .B(_0602_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2003_ (.A1(_1074_),
    .A2(_0976_),
    .A3(_1076_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2004_ (.I(_0974_),
    .Z(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2005_ (.I(_0822_),
    .Z(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2006_ (.A1(_1078_),
    .A2(_0889_),
    .B(_1079_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2007_ (.A1(_0887_),
    .A2(_1049_),
    .B1(_1077_),
    .B2(_1080_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2008_ (.A1(_1073_),
    .A2(_1081_),
    .ZN(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2009_ (.A1(_1034_),
    .A2(_1041_),
    .B(_0789_),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2010_ (.A1(_0967_),
    .A2(_0631_),
    .A3(_0847_),
    .ZN(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2011_ (.A1(_0820_),
    .A2(_0916_),
    .A3(_0969_),
    .ZN(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2012_ (.A1(_0739_),
    .A2(_0854_),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2013_ (.A1(_0967_),
    .A2(_0732_),
    .A3(_1086_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2014_ (.A1(_1085_),
    .A2(_1087_),
    .B(_1084_),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2015_ (.A1(_1084_),
    .A2(_1085_),
    .B(_1088_),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2016_ (.I(_0812_),
    .Z(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2017_ (.A1(_1090_),
    .A2(_0754_),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2018_ (.A1(_0771_),
    .A2(_1089_),
    .B1(_1091_),
    .B2(_0500_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2019_ (.A1(_1083_),
    .A2(_1092_),
    .Z(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2020_ (.I(_1044_),
    .Z(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2021_ (.A1(_0666_),
    .A2(_0710_),
    .B(_1025_),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2022_ (.A1(_0666_),
    .A2(_0710_),
    .B(_1095_),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2023_ (.A1(_0807_),
    .A2(_0969_),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2024_ (.A1(_0844_),
    .A2(_0971_),
    .A3(_1075_),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2025_ (.A1(_0893_),
    .A2(_1097_),
    .B(_1098_),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _2026_ (.A1(_0820_),
    .A2(_0782_),
    .A3(_0989_),
    .B1(_1097_),
    .B2(_1098_),
    .B3(_0893_),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2027_ (.A1(_1029_),
    .A2(net46),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2028_ (.A1(_1079_),
    .A2(_1096_),
    .B1(_1099_),
    .B2(_1101_),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2029_ (.A1(_1056_),
    .A2(_1102_),
    .Z(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2030_ (.I(_1044_),
    .Z(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2031_ (.A1(_1104_),
    .A2(_1057_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2032_ (.A1(_1094_),
    .A2(_1103_),
    .B(_1105_),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2033_ (.A1(_0925_),
    .A2(_1093_),
    .B(_1106_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2034_ (.A1(_1083_),
    .A2(_1092_),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2035_ (.A1(_0997_),
    .A2(_1059_),
    .B(_0863_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2036_ (.I0(_1109_),
    .I1(_1103_),
    .S(_0942_),
    .Z(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2037_ (.A1(_0730_),
    .A2(_1108_),
    .A3(_1110_),
    .B(_0672_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2038_ (.A1(_1082_),
    .A2(_1107_),
    .A3(_1111_),
    .Z(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2039_ (.A1(_1107_),
    .A2(_1111_),
    .B(_1082_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2040_ (.A1(_1112_),
    .A2(_1113_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2041_ (.A1(_1071_),
    .A2(_1114_),
    .Z(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2042_ (.A1(_1015_),
    .A2(_1014_),
    .A3(_1017_),
    .A4(_1067_),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2043_ (.A1(_1020_),
    .A2(_1021_),
    .B(_1066_),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2044_ (.A1(_1020_),
    .A2(_1021_),
    .A3(_1066_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2045_ (.A1(_1068_),
    .A2(_1117_),
    .B(_1118_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2046_ (.A1(_1116_),
    .A2(_1119_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2047_ (.A1(_1115_),
    .A2(_1120_),
    .Z(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2048_ (.I(_1121_),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2049_ (.I(_0925_),
    .Z(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2050_ (.A1(_1122_),
    .A2(_1093_),
    .A3(_1106_),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2051_ (.A1(_0960_),
    .A2(_1082_),
    .A3(_1107_),
    .B(_1123_),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2052_ (.I(_1079_),
    .Z(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2053_ (.I(_0808_),
    .Z(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2054_ (.A1(_1038_),
    .A2(_0968_),
    .ZN(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2055_ (.A1(_1126_),
    .A2(_1127_),
    .B(_1087_),
    .C(_0874_),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2056_ (.I(_1079_),
    .Z(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2057_ (.A1(_1129_),
    .A2(_0969_),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2058_ (.I(_0604_),
    .Z(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2059_ (.A1(_1125_),
    .A2(_1128_),
    .B(_1130_),
    .C(_1131_),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2060_ (.A1(_1073_),
    .A2(_1132_),
    .Z(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2061_ (.I(_1090_),
    .Z(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2062_ (.A1(_0826_),
    .A2(_1023_),
    .B1(_0911_),
    .B2(_1134_),
    .C(_0974_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2063_ (.A1(_0660_),
    .A2(_0714_),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2064_ (.A1(_0809_),
    .A2(_1136_),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2065_ (.A1(_0928_),
    .A2(_1137_),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2066_ (.A1(_0936_),
    .A2(_1138_),
    .B(_1074_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2067_ (.A1(_0718_),
    .A2(_1003_),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _2068_ (.A1(_1129_),
    .A2(_1135_),
    .A3(_1139_),
    .B1(_0875_),
    .B2(_1140_),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2069_ (.A1(_1109_),
    .A2(_1141_),
    .Z(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2070_ (.A1(_0618_),
    .A2(_1141_),
    .B(_1094_),
    .ZN(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2071_ (.I(_1083_),
    .Z(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2072_ (.A1(_1086_),
    .A2(_0847_),
    .A3(_1137_),
    .ZN(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2073_ (.A1(_0867_),
    .A2(_0849_),
    .B(_1027_),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _2074_ (.A1(_1078_),
    .A2(_1145_),
    .B(_1146_),
    .C(_0771_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2075_ (.A1(_1144_),
    .A2(_1147_),
    .Z(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _2076_ (.A1(_1094_),
    .A2(_0998_),
    .Z(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2077_ (.A1(_1142_),
    .A2(_1143_),
    .B1(_1148_),
    .B2(_0925_),
    .C(_1149_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2078_ (.A1(_1142_),
    .A2(_1143_),
    .B(_1149_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2079_ (.A1(_1144_),
    .A2(_1147_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2080_ (.A1(_0731_),
    .A2(_1151_),
    .A3(_1152_),
    .B(_0672_),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2081_ (.A1(_1133_),
    .A2(_1150_),
    .A3(_1153_),
    .Z(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2082_ (.A1(_1150_),
    .A2(_1153_),
    .B(_1133_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2083_ (.A1(_1124_),
    .A2(_1154_),
    .A3(_1155_),
    .Z(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2084_ (.A1(_1154_),
    .A2(_1155_),
    .B(_1124_),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2085_ (.A1(_1156_),
    .A2(_1157_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2086_ (.A1(_1071_),
    .A2(_1112_),
    .A3(_1113_),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2087_ (.A1(_1115_),
    .A2(_1120_),
    .B(_1159_),
    .ZN(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2088_ (.A1(_1158_),
    .A2(_1160_),
    .Z(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2089_ (.I(_1161_),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2090_ (.I(_1157_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2091_ (.A1(_1124_),
    .A2(_1154_),
    .A3(_1155_),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2092_ (.A1(_1159_),
    .A2(_1163_),
    .ZN(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2093_ (.A1(_1162_),
    .A2(_1164_),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2094_ (.A1(_1071_),
    .A2(_1114_),
    .ZN(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2095_ (.A1(_1116_),
    .A2(_1119_),
    .B(_1158_),
    .C(_1166_),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2096_ (.A1(_0731_),
    .A2(_1151_),
    .A3(_1152_),
    .B(_1154_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2097_ (.A1(_0826_),
    .A2(_1023_),
    .B(_0801_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2098_ (.A1(_1090_),
    .A2(_1025_),
    .A3(_0932_),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2099_ (.A1(_0967_),
    .A2(_0813_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2100_ (.A1(_1090_),
    .A2(_0975_),
    .B1(_1171_),
    .B2(_0927_),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2101_ (.A1(_0928_),
    .A2(_1170_),
    .B1(_1172_),
    .B2(_0808_),
    .C(_1029_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _2102_ (.A1(_1074_),
    .A2(_0646_),
    .A3(_0933_),
    .B1(_1169_),
    .B2(_1173_),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2103_ (.A1(_0863_),
    .A2(_1174_),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2104_ (.A1(_1057_),
    .A2(_1174_),
    .B(_1175_),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2105_ (.A1(_1104_),
    .A2(_0998_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _2106_ (.A1(_1104_),
    .A2(_1176_),
    .B(_1177_),
    .C(_0670_),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2107_ (.I(_0804_),
    .Z(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2108_ (.A1(_0689_),
    .A2(_1023_),
    .ZN(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2109_ (.A1(_1027_),
    .A2(_1180_),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2110_ (.A1(_0808_),
    .A2(_1137_),
    .B(_1029_),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _2111_ (.A1(_0974_),
    .A2(_1051_),
    .B(_1181_),
    .C(_1182_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2112_ (.A1(_1001_),
    .A2(_1034_),
    .A3(_1041_),
    .ZN(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2113_ (.A1(_1179_),
    .A2(_1184_),
    .B(_1183_),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2114_ (.A1(_1179_),
    .A2(_1183_),
    .B(_1185_),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2115_ (.A1(_0730_),
    .A2(_1186_),
    .ZN(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2116_ (.A1(_1178_),
    .A2(_1187_),
    .Z(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2117_ (.A1(_0562_),
    .A2(_0624_),
    .A3(_0604_),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2118_ (.A1(_0809_),
    .A2(_0970_),
    .ZN(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2119_ (.A1(_1075_),
    .A2(_0855_),
    .B(_0602_),
    .ZN(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2120_ (.A1(_1078_),
    .A2(_1190_),
    .A3(_1191_),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2121_ (.A1(_1072_),
    .A2(_1192_),
    .B(_1189_),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2122_ (.I0(_1189_),
    .I1(_1193_),
    .S(_0619_),
    .Z(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2123_ (.I(_1194_),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2124_ (.A1(_1188_),
    .A2(_1195_),
    .Z(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2125_ (.A1(_1168_),
    .A2(_1196_),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2126_ (.A1(_1165_),
    .A2(_1167_),
    .B(_1197_),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2127_ (.A1(_1197_),
    .A2(_1165_),
    .A3(_1167_),
    .Z(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2128_ (.A1(_1198_),
    .A2(_1199_),
    .ZN(net28));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2129_ (.A1(_0731_),
    .A2(_1178_),
    .A3(_1186_),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2130_ (.A1(_1188_),
    .A2(_1195_),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2131_ (.I(_1125_),
    .Z(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2132_ (.A1(_0889_),
    .A2(_0511_),
    .ZN(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2133_ (.I(_1203_),
    .ZN(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2134_ (.A1(_1202_),
    .A2(_1204_),
    .B(_0624_),
    .C(_1131_),
    .ZN(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2135_ (.A1(_1031_),
    .A2(_1205_),
    .ZN(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2136_ (.A1(_1073_),
    .A2(_1205_),
    .B(_1206_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2137_ (.A1(_0660_),
    .A2(_0663_),
    .B(_0975_),
    .C(_1134_),
    .ZN(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2138_ (.A1(_1126_),
    .A2(_0689_),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2139_ (.A1(_1126_),
    .A2(_1051_),
    .B1(_1208_),
    .B2(_1209_),
    .C(_1129_),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2140_ (.A1(_1125_),
    .A2(_1192_),
    .B(_1210_),
    .ZN(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2141_ (.A1(_1109_),
    .A2(_1211_),
    .ZN(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2142_ (.A1(_0618_),
    .A2(_1211_),
    .B(_1212_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2143_ (.I(_0671_),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2144_ (.A1(_1094_),
    .A2(_1213_),
    .B(_1177_),
    .C(_0022_),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2145_ (.A1(_1204_),
    .A2(_1136_),
    .B(_1078_),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2146_ (.A1(_1182_),
    .A2(_1215_),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2147_ (.A1(_1144_),
    .A2(_1216_),
    .ZN(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2148_ (.A1(_1179_),
    .A2(_1216_),
    .B(_1217_),
    .C(_1122_),
    .ZN(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2149_ (.A1(_1214_),
    .A2(_1218_),
    .Z(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2150_ (.A1(_1207_),
    .A2(_1219_),
    .Z(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2151_ (.A1(_1200_),
    .A2(_1201_),
    .B(_1220_),
    .ZN(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2152_ (.A1(_1200_),
    .A2(_1201_),
    .A3(_1220_),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2153_ (.I(_1222_),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2154_ (.A1(_1221_),
    .A2(_1223_),
    .ZN(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2155_ (.A1(_1168_),
    .A2(_1196_),
    .B(_1198_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2156_ (.A1(_1224_),
    .A2(_1225_),
    .Z(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2157_ (.I(_1226_),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2158_ (.I(_1074_),
    .Z(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2159_ (.A1(_1126_),
    .A2(_0914_),
    .A3(_0712_),
    .B(_1129_),
    .ZN(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2160_ (.A1(_1125_),
    .A2(_1227_),
    .A3(_1039_),
    .B(_1228_),
    .ZN(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2161_ (.A1(_1104_),
    .A2(_1057_),
    .Z(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2162_ (.A1(_1229_),
    .A2(_1230_),
    .Z(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2163_ (.A1(_0022_),
    .A2(_1231_),
    .ZN(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2164_ (.A1(_1227_),
    .A2(_0734_),
    .B(_1182_),
    .ZN(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2165_ (.A1(_1144_),
    .A2(_1233_),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _2166_ (.A1(_1179_),
    .A2(_1233_),
    .B(_1234_),
    .C(_1122_),
    .ZN(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2167_ (.A1(_1232_),
    .A2(_1235_),
    .Z(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2168_ (.A1(_1232_),
    .A2(_1235_),
    .ZN(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2169_ (.A1(_1236_),
    .A2(_1237_),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2170_ (.A1(_1131_),
    .A2(_1073_),
    .ZN(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2171_ (.I(_0624_),
    .ZN(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2172_ (.A1(_1031_),
    .A2(_1131_),
    .B(_1239_),
    .C(_1240_),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2173_ (.I(_1241_),
    .Z(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2174_ (.A1(_1238_),
    .A2(_1242_),
    .Z(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2175_ (.A1(_1238_),
    .A2(_1242_),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2176_ (.A1(_1243_),
    .A2(_1244_),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2177_ (.A1(_1214_),
    .A2(_1218_),
    .ZN(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2178_ (.A1(_1207_),
    .A2(_1219_),
    .B(_1246_),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _2179_ (.A1(_1245_),
    .A2(_1247_),
    .ZN(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2180_ (.A1(_1168_),
    .A2(_1196_),
    .ZN(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2181_ (.A1(_1249_),
    .A2(_1221_),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2182_ (.A1(_1198_),
    .A2(_1250_),
    .ZN(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2183_ (.A1(_1222_),
    .A2(_1251_),
    .ZN(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2184_ (.A1(_1248_),
    .A2(_1252_),
    .ZN(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2185_ (.I(_1253_),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2186_ (.A1(_1134_),
    .A2(_0968_),
    .B(_1227_),
    .ZN(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2187_ (.A1(_1134_),
    .A2(_0754_),
    .B1(_1254_),
    .B2(_1202_),
    .ZN(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2188_ (.A1(_0618_),
    .A2(_1255_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2189_ (.A1(_1109_),
    .A2(_1255_),
    .B(_1256_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2190_ (.A1(_0942_),
    .A2(_1257_),
    .B(_1149_),
    .C(_0960_),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2191_ (.A1(_1235_),
    .A2(_1241_),
    .A3(_1259_),
    .ZN(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2192_ (.A1(_1236_),
    .A2(_1243_),
    .B(_1260_),
    .ZN(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2193_ (.A1(_1236_),
    .A2(_1243_),
    .A3(_1260_),
    .Z(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2194_ (.A1(_1261_),
    .A2(_1262_),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2195_ (.A1(_1222_),
    .A2(_1248_),
    .A3(_1251_),
    .B1(_1245_),
    .B2(_1247_),
    .ZN(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2196_ (.A1(_1263_),
    .A2(_1264_),
    .Z(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2197_ (.I(_1265_),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2198_ (.A1(_1242_),
    .A2(_1259_),
    .ZN(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2199_ (.A1(_1242_),
    .A2(_1259_),
    .B(_1235_),
    .ZN(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2200_ (.A1(_1266_),
    .A2(_1267_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2201_ (.I(_1263_),
    .ZN(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2202_ (.A1(_1222_),
    .A2(_1248_),
    .A3(_1251_),
    .A4(_1270_),
    .ZN(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2203_ (.A1(_1245_),
    .A2(_1247_),
    .ZN(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2204_ (.A1(_1236_),
    .A2(_1243_),
    .A3(_1260_),
    .ZN(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2205_ (.A1(_1272_),
    .A2(_1273_),
    .B(_1261_),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2206_ (.I(_1274_),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _2207_ (.A1(_1269_),
    .A2(_1271_),
    .A3(_1275_),
    .B1(_1230_),
    .B2(_0960_),
    .ZN(net20));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2208_ (.A1(_0751_),
    .A2(_0836_),
    .Z(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2209_ (.I(_1276_),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2210_ (.I(_0135_),
    .Z(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2211_ (.I(_1278_),
    .Z(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2212_ (.I(_1408_),
    .Z(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2213_ (.I(_1280_),
    .Z(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2214_ (.I(net55),
    .Z(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2215_ (.I(_1354_),
    .Z(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2216_ (.A1(_1282_),
    .A2(_1283_),
    .B(_0091_),
    .ZN(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2217_ (.I(_1284_),
    .Z(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2218_ (.I(_1321_),
    .Z(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2219_ (.I(_1286_),
    .Z(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2220_ (.I(_1430_),
    .Z(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2221_ (.I(_1289_),
    .Z(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2222_ (.A1(_0157_),
    .A2(_0047_),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2223_ (.I(_0091_),
    .Z(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2224_ (.A1(_1287_),
    .A2(_1290_),
    .B(_1291_),
    .C(_1292_),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2225_ (.I(_1343_),
    .Z(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2226_ (.I(_1354_),
    .Z(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2227_ (.I(_1295_),
    .Z(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2228_ (.A1(_1294_),
    .A2(_1296_),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2229_ (.I(_1268_),
    .Z(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2230_ (.I(_0058_),
    .Z(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2231_ (.A1(_1298_),
    .A2(_1300_),
    .B(_1284_),
    .ZN(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2232_ (.A1(_0157_),
    .A2(_0047_),
    .ZN(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2233_ (.I(_1302_),
    .Z(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _2234_ (.A1(_1281_),
    .A2(_1285_),
    .B1(_1293_),
    .B2(_1297_),
    .C1(_1301_),
    .C2(_1303_),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2235_ (.I(_1268_),
    .Z(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2236_ (.I(_1305_),
    .Z(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2237_ (.I(_1283_),
    .Z(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2238_ (.I(_0091_),
    .Z(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2239_ (.A1(_1306_),
    .A2(_1307_),
    .B(_1308_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2240_ (.I(_1289_),
    .Z(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2241_ (.A1(_1258_),
    .A2(_1321_),
    .Z(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2242_ (.I(_1312_),
    .Z(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2243_ (.I(_0069_),
    .Z(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2244_ (.A1(_1311_),
    .A2(_1313_),
    .B(_1314_),
    .C(_1310_),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2245_ (.I(_0200_),
    .Z(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2246_ (.I(_0124_),
    .Z(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2247_ (.A1(_1316_),
    .A2(_1317_),
    .ZN(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2248_ (.A1(_1309_),
    .A2(_1315_),
    .B(_1318_),
    .ZN(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2249_ (.A1(_1279_),
    .A2(_1304_),
    .B(_1319_),
    .C(_0146_),
    .ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2250_ (.I(_1320_),
    .Z(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2251_ (.I(\p_shaping_I.counter[1] ),
    .ZN(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2252_ (.I(_1323_),
    .Z(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _2253_ (.A1(net31),
    .A2(net30),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2254_ (.I(_0178_),
    .Z(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2255_ (.A1(_1441_),
    .A2(_1325_),
    .B(_0102_),
    .C(_1326_),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2256_ (.A1(_1300_),
    .A2(_1291_),
    .B(_1299_),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _2257_ (.A1(_0211_),
    .A2(_1408_),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2258_ (.A1(_1327_),
    .A2(_1328_),
    .B(_1329_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2259_ (.I(_0178_),
    .Z(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2260_ (.A1(_1331_),
    .A2(_1291_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2261_ (.A1(_1280_),
    .A2(_1333_),
    .B(_0211_),
    .ZN(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2262_ (.I(_1258_),
    .Z(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2263_ (.I(_1321_),
    .Z(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _2264_ (.A1(_1335_),
    .A2(_1336_),
    .Z(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2265_ (.A1(_1335_),
    .A2(_1282_),
    .B(_1365_),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2266_ (.A1(_1331_),
    .A2(_1338_),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _2267_ (.A1(_1305_),
    .A2(_1289_),
    .B(_1336_),
    .ZN(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2268_ (.A1(_0211_),
    .A2(_0124_),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2269_ (.A1(_1337_),
    .A2(_1339_),
    .B1(_1340_),
    .B2(_1308_),
    .C(_1341_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2270_ (.A1(_1330_),
    .A2(_1334_),
    .A3(_1342_),
    .Z(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2271_ (.I(_1344_),
    .Z(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2272_ (.I(_0124_),
    .Z(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _2273_ (.A1(_0036_),
    .A2(_0047_),
    .A3(net33),
    .A4(_0058_),
    .Z(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2274_ (.A1(_1346_),
    .A2(_1347_),
    .B(_1316_),
    .ZN(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2275_ (.I(_1308_),
    .Z(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2276_ (.A1(_0036_),
    .A2(_1430_),
    .ZN(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2277_ (.I(_1350_),
    .Z(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2278_ (.I0(_1349_),
    .I1(_1309_),
    .S(_1351_),
    .Z(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2279_ (.I(_0036_),
    .Z(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2280_ (.I(_1353_),
    .Z(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2281_ (.I(_1307_),
    .Z(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2282_ (.A1(_1355_),
    .A2(_1294_),
    .B(_1356_),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2283_ (.I(_1289_),
    .Z(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2284_ (.I(_1358_),
    .Z(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2285_ (.A1(_1353_),
    .A2(_1286_),
    .Z(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2286_ (.I(_1360_),
    .Z(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2287_ (.I(_1288_),
    .Z(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2288_ (.I(_1362_),
    .Z(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2289_ (.A1(_1359_),
    .A2(_1361_),
    .B(_1363_),
    .ZN(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2290_ (.I(_0178_),
    .Z(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2291_ (.I(_1366_),
    .Z(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2292_ (.I(_1325_),
    .Z(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _2293_ (.A1(_1335_),
    .A2(_1365_),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2294_ (.A1(_1367_),
    .A2(_1368_),
    .A3(_1369_),
    .ZN(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2295_ (.I(_1408_),
    .Z(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2296_ (.I(_1371_),
    .Z(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2297_ (.A1(_1357_),
    .A2(_1364_),
    .B(_1370_),
    .C(_1372_),
    .ZN(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2298_ (.I(_1362_),
    .Z(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2299_ (.I(_1337_),
    .Z(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2300_ (.A1(_1374_),
    .A2(_1375_),
    .A3(_1369_),
    .ZN(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2301_ (.I(_1346_),
    .Z(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2302_ (.I(_1282_),
    .Z(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2303_ (.A1(_1379_),
    .A2(_1366_),
    .A3(_1300_),
    .ZN(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2304_ (.A1(_1378_),
    .A2(_1380_),
    .Z(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2305_ (.I(_0135_),
    .Z(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2306_ (.I(_1382_),
    .Z(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2307_ (.A1(_1377_),
    .A2(_1381_),
    .B(_1383_),
    .ZN(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2308_ (.A1(_1348_),
    .A2(_1352_),
    .B1(_1373_),
    .B2(_1384_),
    .ZN(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2309_ (.I(_1385_),
    .Z(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2310_ (.A1(_1324_),
    .A2(_1345_),
    .B(_1386_),
    .ZN(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2311_ (.I(\p_shaping_I.counter[1] ),
    .Z(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2312_ (.A1(_1389_),
    .A2(\p_shaping_I.counter[0] ),
    .ZN(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2313_ (.I(_1390_),
    .ZN(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2314_ (.A1(_1324_),
    .A2(_1386_),
    .A3(_1345_),
    .Z(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2315_ (.A1(_1388_),
    .A2(_1391_),
    .A3(_1392_),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2316_ (.A1(_1322_),
    .A2(_1393_),
    .Z(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2317_ (.I(_1394_),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2318_ (.A1(_1322_),
    .A2(_1393_),
    .Z(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2319_ (.A1(_1392_),
    .A2(_1395_),
    .Z(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2320_ (.I(_1382_),
    .Z(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2321_ (.I(_1286_),
    .Z(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2322_ (.A1(_1277_),
    .A2(_1399_),
    .ZN(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2323_ (.I(_1283_),
    .Z(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2324_ (.I(_1305_),
    .Z(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _2325_ (.A1(_1379_),
    .A2(_1401_),
    .B(_1402_),
    .ZN(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2326_ (.I(_1346_),
    .Z(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _2327_ (.I0(_1314_),
    .I1(_0113_),
    .I2(_1400_),
    .I3(_1403_),
    .S0(_1404_),
    .S1(_1363_),
    .Z(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2328_ (.I(_1404_),
    .Z(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2329_ (.I(_1338_),
    .Z(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2330_ (.A1(_1296_),
    .A2(_1313_),
    .B(_1407_),
    .C(_1349_),
    .ZN(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2331_ (.A1(_1406_),
    .A2(_1301_),
    .A3(_1409_),
    .B(_1279_),
    .ZN(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2332_ (.A1(_1398_),
    .A2(_1405_),
    .B(_1410_),
    .ZN(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2333_ (.A1(\p_shaping_I.bit_in ),
    .A2(_1322_),
    .ZN(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2334_ (.A1(_1411_),
    .A2(_1412_),
    .ZN(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2335_ (.A1(\p_shaping_I.bit_in_2 ),
    .A2(_1330_),
    .A3(_1334_),
    .A4(_1342_),
    .ZN(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _2336_ (.A1(_1353_),
    .A2(_1343_),
    .B(_1441_),
    .ZN(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2337_ (.A1(_1298_),
    .A2(_1326_),
    .A3(_1300_),
    .ZN(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2338_ (.I(_1336_),
    .Z(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2339_ (.A1(_1292_),
    .A2(_1415_),
    .B1(_1416_),
    .B2(_1417_),
    .ZN(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2340_ (.A1(_1376_),
    .A2(_1312_),
    .B(_1331_),
    .ZN(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2341_ (.A1(_1301_),
    .A2(_1420_),
    .B(_1280_),
    .ZN(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2342_ (.I(_0189_),
    .Z(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2343_ (.A1(_1422_),
    .A2(_1325_),
    .ZN(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2344_ (.A1(_1278_),
    .A2(_1423_),
    .ZN(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2345_ (.A1(_1348_),
    .A2(_1418_),
    .B1(_1421_),
    .B2(_1424_),
    .ZN(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2346_ (.I(_1425_),
    .Z(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2347_ (.A1(_1414_),
    .A2(_1426_),
    .Z(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2348_ (.I(_0607_),
    .Z(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2349_ (.I(_1347_),
    .Z(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2350_ (.A1(_1317_),
    .A2(_1429_),
    .ZN(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2351_ (.A1(_1278_),
    .A2(_1431_),
    .ZN(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2352_ (.I(_1295_),
    .Z(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2353_ (.A1(_1306_),
    .A2(_1362_),
    .A3(_1433_),
    .ZN(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2354_ (.A1(_1309_),
    .A2(_1351_),
    .B(_1434_),
    .ZN(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2355_ (.A1(_1306_),
    .A2(_1287_),
    .B(_1290_),
    .ZN(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2356_ (.A1(_1401_),
    .A2(_1303_),
    .B(_1308_),
    .ZN(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2357_ (.I(_1288_),
    .Z(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2358_ (.A1(_1353_),
    .A2(_1295_),
    .Z(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2359_ (.A1(_1438_),
    .A2(_1439_),
    .ZN(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2360_ (.A1(_1436_),
    .A2(_1437_),
    .B1(_1440_),
    .B2(_1368_),
    .C(_1404_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2361_ (.I(_1291_),
    .Z(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2362_ (.A1(_1292_),
    .A2(_0027_),
    .A3(_1439_),
    .B(_1380_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2363_ (.A1(_1371_),
    .A2(_0028_),
    .B(_1316_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2364_ (.A1(_1432_),
    .A2(_1435_),
    .B1(_0026_),
    .B2(_0029_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2365_ (.I(_1430_),
    .Z(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _2366_ (.A1(_0031_),
    .A2(_1368_),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2367_ (.A1(_1433_),
    .A2(_1337_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2368_ (.I(_1438_),
    .Z(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2369_ (.A1(_0032_),
    .A2(_0033_),
    .B(_0034_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2370_ (.A1(_1402_),
    .A2(_1417_),
    .A3(_1307_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2371_ (.A1(_1372_),
    .A2(_0032_),
    .A3(_0037_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2372_ (.I(_1326_),
    .Z(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2373_ (.A1(_0039_),
    .A2(_0113_),
    .B(_1317_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _2374_ (.A1(_0035_),
    .A2(_0038_),
    .B(_1398_),
    .C(_0040_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2375_ (.A1(_1311_),
    .A2(_1337_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2376_ (.A1(_1305_),
    .A2(_1336_),
    .B(_1283_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2377_ (.I(_0043_),
    .Z(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2378_ (.A1(_0042_),
    .A2(_0044_),
    .B(_1349_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2379_ (.I(_1378_),
    .Z(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2380_ (.A1(_1282_),
    .A2(_0058_),
    .Z(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2381_ (.A1(_1402_),
    .A2(_1417_),
    .A3(_1401_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2382_ (.A1(_0046_),
    .A2(_0048_),
    .A3(_0049_),
    .Z(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2383_ (.I(_1299_),
    .Z(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2384_ (.I(_0051_),
    .Z(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2385_ (.A1(_0052_),
    .A2(_1314_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2386_ (.I(_1355_),
    .Z(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2387_ (.I(_1367_),
    .Z(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2388_ (.A1(_0054_),
    .A2(_1359_),
    .B(_0055_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2389_ (.A1(_0053_),
    .A2(_0056_),
    .B(_0046_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2390_ (.I(_1316_),
    .Z(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _2391_ (.A1(_0045_),
    .A2(_0050_),
    .B(_0057_),
    .C(_0059_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2392_ (.A1(_1428_),
    .A2(_0030_),
    .A3(_0041_),
    .A4(_0060_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2393_ (.I(\p_shaping_I.bit_in_1 ),
    .Z(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2394_ (.I(_0062_),
    .Z(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2395_ (.A1(_1296_),
    .A2(_1313_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2396_ (.A1(_1311_),
    .A2(_0027_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2397_ (.A1(_0064_),
    .A2(_0065_),
    .B(_1367_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2398_ (.A1(_1371_),
    .A2(_0032_),
    .A3(_0037_),
    .Z(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2399_ (.A1(_1382_),
    .A2(_0040_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2400_ (.A1(_0066_),
    .A2(_0067_),
    .B(_0068_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2401_ (.A1(_1433_),
    .A2(_0027_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2402_ (.I(_1332_),
    .Z(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2403_ (.A1(_1355_),
    .A2(_0072_),
    .B(_1290_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2404_ (.A1(_0071_),
    .A2(_0073_),
    .B(_0034_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2405_ (.A1(_1404_),
    .A2(_0048_),
    .A3(_0049_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2406_ (.A1(_1335_),
    .A2(_1286_),
    .A3(_1295_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2407_ (.A1(_0039_),
    .A2(_0076_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2408_ (.A1(_1402_),
    .A2(_1307_),
    .B(_1362_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2409_ (.A1(_0077_),
    .A2(_0078_),
    .B(_1371_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2410_ (.A1(_0074_),
    .A2(_0075_),
    .B(_0079_),
    .C(_1382_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2411_ (.A1(_0063_),
    .A2(_1386_),
    .B1(_0070_),
    .B2(_0081_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2412_ (.A1(_1323_),
    .A2(_1427_),
    .B(_0061_),
    .C(_0082_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2413_ (.A1(_1428_),
    .A2(_0030_),
    .B1(_0041_),
    .B2(_0060_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2414_ (.A1(_0062_),
    .A2(_1386_),
    .A3(_0070_),
    .A4(_0081_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2415_ (.A1(_1414_),
    .A2(_1426_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2416_ (.A1(_0084_),
    .A2(_0085_),
    .B(_0086_),
    .C(_1389_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2417_ (.A1(_1391_),
    .A2(_0083_),
    .A3(_0087_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2418_ (.A1(_1413_),
    .A2(_0088_),
    .Z(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2419_ (.A1(_1396_),
    .A2(_0089_),
    .Z(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2420_ (.I(_1413_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2421_ (.A1(_0092_),
    .A2(_0088_),
    .B(_0087_),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2422_ (.I(\p_shaping_I.bit_in ),
    .Z(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2423_ (.A1(_1322_),
    .A2(_1411_),
    .B(_0094_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2424_ (.A1(_1278_),
    .A2(_1280_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2425_ (.A1(_1356_),
    .A2(_1303_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2426_ (.A1(_0055_),
    .A2(_0097_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2427_ (.A1(_0096_),
    .A2(_0032_),
    .A3(_0098_),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2428_ (.I(_1294_),
    .Z(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2429_ (.I(_1331_),
    .Z(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2430_ (.A1(_0101_),
    .A2(_1340_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2431_ (.A1(_0100_),
    .A2(_0078_),
    .B(_0103_),
    .C(_1318_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2432_ (.A1(_1376_),
    .A2(_1302_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2433_ (.I(_0157_),
    .Z(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _2434_ (.A1(_0106_),
    .A2(_1343_),
    .A3(_1441_),
    .B(_1438_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2435_ (.A1(_0135_),
    .A2(_1346_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2436_ (.I(_0108_),
    .Z(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2437_ (.A1(_0105_),
    .A2(_0107_),
    .B(_0077_),
    .C(_0109_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2438_ (.A1(_0099_),
    .A2(_0104_),
    .A3(_0110_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2439_ (.A1(_0095_),
    .A2(_0111_),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2440_ (.I(_1391_),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2441_ (.I(_1324_),
    .Z(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2442_ (.I(\p_shaping_I.bit_in_2 ),
    .Z(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2443_ (.A1(_1345_),
    .A2(_1426_),
    .B(_0116_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2444_ (.A1(_1314_),
    .A2(_1338_),
    .B1(_1415_),
    .B2(_0101_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2445_ (.A1(_0051_),
    .A2(_0105_),
    .B(_1341_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2446_ (.A1(_1298_),
    .A2(_1379_),
    .B(_1438_),
    .C(_0031_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2447_ (.I(_1419_),
    .Z(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2448_ (.A1(_1380_),
    .A2(_0120_),
    .B(_0121_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2449_ (.A1(_1298_),
    .A2(_1379_),
    .A3(_1366_),
    .A4(_1376_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2450_ (.A1(_1326_),
    .A2(_0048_),
    .Z(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2451_ (.A1(_0108_),
    .A2(_1415_),
    .A3(_0123_),
    .A4(_0125_),
    .Z(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2452_ (.A1(_0118_),
    .A2(_0119_),
    .B(_0122_),
    .C(_0126_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2453_ (.A1(_0117_),
    .A2(_0127_),
    .Z(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2454_ (.A1(_1367_),
    .A2(_1403_),
    .B(_1420_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2455_ (.I(_1317_),
    .Z(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2456_ (.A1(_0106_),
    .A2(_1366_),
    .Z(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2457_ (.A1(_0072_),
    .A2(_1296_),
    .A3(_0131_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2458_ (.A1(_0130_),
    .A2(_0132_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2459_ (.A1(_1406_),
    .A2(_0129_),
    .B(_0133_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2460_ (.A1(_1417_),
    .A2(_1358_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2461_ (.A1(_1333_),
    .A2(_0136_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2462_ (.A1(_0072_),
    .A2(_1292_),
    .A3(_1369_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2463_ (.A1(_0096_),
    .A2(_0138_),
    .Z(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2464_ (.I(_0108_),
    .Z(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2465_ (.A1(_0072_),
    .A2(_0031_),
    .B(_0106_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2466_ (.A1(_1306_),
    .A2(_1433_),
    .B(_1287_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _2467_ (.A1(_0034_),
    .A2(_0141_),
    .B1(_0107_),
    .B2(_0142_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2468_ (.A1(_0140_),
    .A2(_0143_),
    .Z(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2469_ (.A1(_1398_),
    .A2(_0134_),
    .B1(_0137_),
    .B2(_0139_),
    .C(_0144_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2470_ (.A1(_0610_),
    .A2(_0613_),
    .Z(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2471_ (.A1(_0254_),
    .A2(_0147_),
    .Z(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2472_ (.I(_0148_),
    .Z(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2473_ (.A1(_1385_),
    .A2(_0041_),
    .A3(_0060_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2474_ (.A1(_0145_),
    .A2(_0149_),
    .B(_0608_),
    .C(_0150_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2475_ (.A1(_0030_),
    .A2(_0070_),
    .A3(_0081_),
    .B(_0606_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2476_ (.I0(_1397_),
    .I1(_0129_),
    .S(_1281_),
    .Z(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2477_ (.A1(_0140_),
    .A2(_0143_),
    .B1(_0137_),
    .B2(_0139_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2478_ (.A1(_0059_),
    .A2(_0153_),
    .B(_0154_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2479_ (.I(_0155_),
    .Z(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2480_ (.A1(_0265_),
    .A2(_0147_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2481_ (.I(_0158_),
    .Z(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2482_ (.A1(_0152_),
    .A2(_0156_),
    .A3(_0159_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2483_ (.A1(_0115_),
    .A2(_0128_),
    .B(_0151_),
    .C(_0160_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2484_ (.I(_0158_),
    .Z(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2485_ (.A1(_0152_),
    .A2(_0156_),
    .A3(_0162_),
    .Z(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2486_ (.A1(_0156_),
    .A2(_0162_),
    .B(_0152_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2487_ (.A1(_0117_),
    .A2(_0127_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2488_ (.I(_1389_),
    .Z(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _2489_ (.A1(_0163_),
    .A2(_0164_),
    .B(_0165_),
    .C(_0166_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2490_ (.A1(_0114_),
    .A2(_0161_),
    .A3(_0167_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2491_ (.A1(_0093_),
    .A2(_0112_),
    .A3(_0169_),
    .Z(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2492_ (.A1(_0090_),
    .A2(_0170_),
    .Z(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2493_ (.I(_0171_),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2494_ (.A1(_0114_),
    .A2(_0112_),
    .A3(_0161_),
    .A4(_0167_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2495_ (.A1(_0167_),
    .A2(_0172_),
    .Z(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2496_ (.I(_0130_),
    .Z(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2497_ (.I(_1285_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2498_ (.I(_1313_),
    .Z(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2499_ (.A1(_0175_),
    .A2(_0176_),
    .B1(_0064_),
    .B2(_1374_),
    .C(_0130_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2500_ (.A1(_0174_),
    .A2(_0132_),
    .B(_0177_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2501_ (.I(_1416_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _2502_ (.A1(_1399_),
    .A2(_1311_),
    .B(_0039_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2503_ (.A1(_1356_),
    .A2(_1375_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2504_ (.A1(_1294_),
    .A2(_0180_),
    .B1(_0181_),
    .B2(_1375_),
    .C(_0182_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2505_ (.I(_1341_),
    .Z(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2506_ (.I(_1349_),
    .Z(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2507_ (.A1(_0185_),
    .A2(_0073_),
    .B(_0103_),
    .C(_0140_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _2508_ (.A1(_0059_),
    .A2(_0179_),
    .B1(_0183_),
    .B2(_0184_),
    .C(_0186_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2509_ (.A1(_1320_),
    .A2(_1411_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2510_ (.A1(_0188_),
    .A2(_0111_),
    .B(_0610_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2511_ (.A1(_0187_),
    .A2(_0190_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2512_ (.I(_0116_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2513_ (.I(_0192_),
    .Z(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2514_ (.A1(_1287_),
    .A2(_1290_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2515_ (.A1(_1401_),
    .A2(_1312_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2516_ (.A1(_0194_),
    .A2(_0195_),
    .B(_0141_),
    .C(_0101_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2517_ (.A1(_0031_),
    .A2(_1368_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2518_ (.A1(_0051_),
    .A2(_1403_),
    .B(_0197_),
    .C(_1387_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2519_ (.A1(_0121_),
    .A2(_0196_),
    .A3(_0198_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2520_ (.A1(_1351_),
    .A2(_0044_),
    .B(_0101_),
    .C(_0027_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2521_ (.A1(_0039_),
    .A2(_1350_),
    .A3(_0043_),
    .Z(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2522_ (.I(_0076_),
    .Z(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2523_ (.A1(_1358_),
    .A2(_1303_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2524_ (.A1(_0106_),
    .A2(_1358_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2525_ (.A1(_0203_),
    .A2(_0204_),
    .B(_1285_),
    .C(_0205_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2526_ (.A1(_1299_),
    .A2(_1369_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _2527_ (.A1(_1387_),
    .A2(_0207_),
    .B(_0108_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2528_ (.A1(_0184_),
    .A2(_0201_),
    .A3(_0202_),
    .B1(_0206_),
    .B2(_0208_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2529_ (.A1(_0199_),
    .A2(_0209_),
    .Z(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2530_ (.A1(_1344_),
    .A2(_1425_),
    .A3(_0127_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2531_ (.A1(_0193_),
    .A2(_0210_),
    .A3(_0212_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2532_ (.A1(_1345_),
    .A2(_1426_),
    .A3(_0127_),
    .Z(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2533_ (.A1(_0199_),
    .A2(_0209_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2534_ (.A1(_0116_),
    .A2(_0214_),
    .B(_0215_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2535_ (.A1(_1389_),
    .A2(_0213_),
    .A3(_0216_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2536_ (.A1(_1310_),
    .A2(_0168_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2537_ (.A1(_1351_),
    .A2(_0044_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2538_ (.A1(_0218_),
    .A2(_0195_),
    .B1(_0219_),
    .B2(_1374_),
    .C(_1378_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2539_ (.I(_0125_),
    .Z(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2540_ (.A1(_1378_),
    .A2(_0103_),
    .A3(_0221_),
    .Z(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2541_ (.A1(_1309_),
    .A2(_0035_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2542_ (.A1(_1383_),
    .A2(_0220_),
    .A3(_0223_),
    .B1(_1432_),
    .B2(_0224_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2543_ (.A1(_0148_),
    .A2(_0225_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2544_ (.A1(_0062_),
    .A2(_0145_),
    .B(_0152_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2545_ (.A1(_0226_),
    .A2(_0227_),
    .Z(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2546_ (.A1(_0217_),
    .A2(_0228_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2547_ (.A1(_1390_),
    .A2(_0229_),
    .Z(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2548_ (.A1(_0191_),
    .A2(_0230_),
    .Z(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2549_ (.I(_1390_),
    .Z(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2550_ (.I(_0166_),
    .Z(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2551_ (.A1(_0234_),
    .A2(_0165_),
    .B(_0164_),
    .C(_0163_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2552_ (.A1(_0160_),
    .A2(_0151_),
    .B(_0128_),
    .C(_0115_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2553_ (.I(_0112_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2554_ (.A1(_0232_),
    .A2(_0235_),
    .A3(_0236_),
    .B(_0237_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2555_ (.A1(_0093_),
    .A2(_0172_),
    .A3(_0238_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2556_ (.A1(_0090_),
    .A2(_0170_),
    .B(_0239_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2557_ (.A1(_0173_),
    .A2(_0231_),
    .A3(_0240_),
    .Z(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2558_ (.I(_0241_),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2559_ (.I(_0191_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2560_ (.A1(_0217_),
    .A2(_0228_),
    .B1(_0230_),
    .B2(_0242_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2561_ (.A1(_0052_),
    .A2(_1439_),
    .A3(_0071_),
    .B(_0221_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2562_ (.A1(_1277_),
    .A2(_1329_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2563_ (.I(_0207_),
    .Z(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2564_ (.A1(_0204_),
    .A2(_0033_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2565_ (.A1(_0055_),
    .A2(_1361_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2566_ (.A1(_0100_),
    .A2(_1359_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2567_ (.A1(_0185_),
    .A2(_0248_),
    .B1(_0249_),
    .B2(_0250_),
    .C(_0121_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2568_ (.A1(_0096_),
    .A2(_0245_),
    .B1(_0246_),
    .B2(_0247_),
    .C(_0251_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2569_ (.A1(_0188_),
    .A2(_0111_),
    .A3(_0187_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2570_ (.A1(_0094_),
    .A2(_0253_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2571_ (.A1(_0252_),
    .A2(_0255_),
    .Z(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2572_ (.A1(_1363_),
    .A2(_1360_),
    .B(_0247_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2573_ (.A1(_0140_),
    .A2(_0257_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2574_ (.A1(_0107_),
    .A2(_0142_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2575_ (.A1(_1355_),
    .A2(_0194_),
    .B(_0136_),
    .C(_0051_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2576_ (.A1(_1279_),
    .A2(_0259_),
    .A3(_0260_),
    .B(_0130_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2577_ (.A1(_1363_),
    .A2(_0195_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2578_ (.A1(_1279_),
    .A2(_1370_),
    .A3(_0262_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2579_ (.A1(_0258_),
    .A2(_0261_),
    .A3(_0263_),
    .Z(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2580_ (.A1(_0210_),
    .A2(_0212_),
    .B(_0264_),
    .C(_0193_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2581_ (.I(_0116_),
    .Z(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2582_ (.A1(_0210_),
    .A2(_0212_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2583_ (.A1(_0258_),
    .A2(_0261_),
    .A3(_0263_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2584_ (.A1(_0267_),
    .A2(_0268_),
    .B(_0269_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2585_ (.A1(_0234_),
    .A2(_0266_),
    .A3(_0270_),
    .Z(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2586_ (.A1(_1400_),
    .A2(_0107_),
    .B(_0181_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2587_ (.A1(_1310_),
    .A2(_1338_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2588_ (.A1(_0138_),
    .A2(_0273_),
    .B(_1281_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2589_ (.A1(_1281_),
    .A2(_0138_),
    .A3(_0273_),
    .Z(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2590_ (.A1(_0272_),
    .A2(_0274_),
    .B(_0275_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2591_ (.A1(_0175_),
    .A2(_0045_),
    .B(_1318_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2592_ (.A1(_1398_),
    .A2(_0276_),
    .B(_0277_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2593_ (.A1(_0155_),
    .A2(_0225_),
    .A3(_0278_),
    .B(_0607_),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2594_ (.I(_0279_),
    .Z(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2595_ (.A1(_0150_),
    .A2(_0156_),
    .A3(_0225_),
    .B(_0608_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2596_ (.I(_1383_),
    .Z(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2597_ (.I(_0282_),
    .Z(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2598_ (.I(_0174_),
    .Z(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2599_ (.I(_0055_),
    .Z(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2600_ (.A1(_1399_),
    .A2(_0205_),
    .B(_0037_),
    .C(_0285_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2601_ (.I(_0174_),
    .Z(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2602_ (.A1(_0168_),
    .A2(_0065_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2603_ (.A1(_0288_),
    .A2(_0289_),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2604_ (.A1(_0284_),
    .A2(_1429_),
    .B1(_0287_),
    .B2(_0290_),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2605_ (.I(_0052_),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2606_ (.I(_1356_),
    .Z(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2607_ (.A1(_0292_),
    .A2(_0293_),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2608_ (.A1(_0054_),
    .A2(_0294_),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2609_ (.A1(_0292_),
    .A2(_0049_),
    .Z(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2610_ (.A1(_0054_),
    .A2(_0100_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _2611_ (.A1(_1329_),
    .A2(_1434_),
    .A3(_0295_),
    .B1(_0296_),
    .B2(_0184_),
    .B3(_0298_),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2612_ (.A1(_0283_),
    .A2(_0291_),
    .B(net45),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2613_ (.A1(_0281_),
    .A2(_0300_),
    .Z(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2614_ (.I0(_0280_),
    .I1(_0301_),
    .S(_0159_),
    .Z(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2615_ (.A1(_0271_),
    .A2(_0302_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2616_ (.A1(_0166_),
    .A2(_0266_),
    .A3(_0270_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2617_ (.A1(_0149_),
    .A2(_0279_),
    .Z(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2618_ (.A1(_0159_),
    .A2(_0301_),
    .B(_0305_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2619_ (.A1(_0304_),
    .A2(_0306_),
    .B(_0232_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2620_ (.A1(_0303_),
    .A2(_0307_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _2621_ (.A1(_0244_),
    .A2(_0256_),
    .A3(_0309_),
    .Z(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2622_ (.A1(_0167_),
    .A2(_0172_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2623_ (.A1(_0242_),
    .A2(_0230_),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2624_ (.A1(_0311_),
    .A2(_0312_),
    .B(_0240_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2625_ (.A1(_0173_),
    .A2(_0231_),
    .B(_0313_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2626_ (.A1(_0310_),
    .A2(_0314_),
    .Z(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2627_ (.I(_0315_),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2628_ (.I(_0256_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2629_ (.A1(_0304_),
    .A2(_0306_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2630_ (.A1(_0316_),
    .A2(_0307_),
    .B(_0317_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2631_ (.A1(_0292_),
    .A2(_0048_),
    .A3(_0049_),
    .B(_0247_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2632_ (.A1(_0288_),
    .A2(_0294_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2633_ (.A1(_0284_),
    .A2(_0320_),
    .B(_0321_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2634_ (.I(_0064_),
    .Z(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2635_ (.I(_1406_),
    .Z(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2636_ (.A1(_0185_),
    .A2(_0293_),
    .B(_0324_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2637_ (.A1(_0323_),
    .A2(_0221_),
    .B(_0325_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2638_ (.A1(_0282_),
    .A2(_1429_),
    .A3(_0326_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2639_ (.A1(_0283_),
    .A2(_0322_),
    .B(_0327_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2640_ (.A1(_0252_),
    .A2(_0253_),
    .Z(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2641_ (.A1(_0094_),
    .A2(_0330_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2642_ (.A1(_0328_),
    .A2(_0331_),
    .Z(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2643_ (.A1(_0210_),
    .A2(_0212_),
    .A3(_0264_),
    .B(_0192_),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2644_ (.A1(_1357_),
    .A2(_1364_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2645_ (.A1(_0109_),
    .A2(_0181_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2646_ (.A1(_0034_),
    .A2(_0203_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2647_ (.A1(_1374_),
    .A2(_1407_),
    .B(_0336_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2648_ (.A1(_0046_),
    .A2(_0337_),
    .B(_1383_),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2649_ (.A1(_0168_),
    .A2(_1377_),
    .B(_1370_),
    .C(_1406_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _2650_ (.A1(_0334_),
    .A2(_0335_),
    .B(_0338_),
    .C(_0339_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2651_ (.A1(_0155_),
    .A2(_0225_),
    .B(_0607_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2652_ (.I(_0278_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2653_ (.A1(_1428_),
    .A2(_0278_),
    .Z(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2654_ (.A1(_0342_),
    .A2(_0343_),
    .B(_0344_),
    .C(_0149_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2655_ (.A1(_0333_),
    .A2(_0341_),
    .B(_1323_),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _2656_ (.A1(_0333_),
    .A2(_0341_),
    .B1(_0345_),
    .B2(_0305_),
    .C(_0346_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2657_ (.A1(_0333_),
    .A2(_0341_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2658_ (.I0(_0608_),
    .I1(_0342_),
    .S(_0343_),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2659_ (.I(_0148_),
    .Z(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2660_ (.A1(_0149_),
    .A2(_0280_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _2661_ (.A1(_1324_),
    .A2(_0348_),
    .B1(_0349_),
    .B2(_0350_),
    .C(_0352_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2662_ (.A1(_1391_),
    .A2(_0347_),
    .A3(_0353_),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2663_ (.A1(_0332_),
    .A2(_0354_),
    .ZN(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2664_ (.A1(_0319_),
    .A2(_0355_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2665_ (.A1(_0316_),
    .A2(_0303_),
    .A3(_0307_),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2666_ (.I(_0114_),
    .Z(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2667_ (.A1(_0271_),
    .A2(_0302_),
    .B(_0025_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2668_ (.A1(_0317_),
    .A2(_0358_),
    .B(_0256_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2669_ (.A1(_0244_),
    .A2(_0357_),
    .A3(_0359_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2670_ (.A1(_0310_),
    .A2(_0314_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2671_ (.A1(_0360_),
    .A2(_0362_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2672_ (.A1(_0356_),
    .A2(_0363_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2673_ (.I(_0364_),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2674_ (.A1(_0332_),
    .A2(_0354_),
    .Z(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2675_ (.A1(_0347_),
    .A2(_0365_),
    .Z(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2676_ (.A1(_0328_),
    .A2(_0330_),
    .B(_0094_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2677_ (.I(_0288_),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2678_ (.I(_1359_),
    .Z(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2679_ (.I(_0285_),
    .Z(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2680_ (.A1(_0369_),
    .A2(_0176_),
    .B(_0113_),
    .C(_0370_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2681_ (.A1(_0368_),
    .A2(_0247_),
    .A3(_0372_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2682_ (.I(_0282_),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2683_ (.I(_0374_),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2684_ (.A1(_0375_),
    .A2(_0325_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2685_ (.A1(_1318_),
    .A2(_0272_),
    .B1(_0373_),
    .B2(_0376_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2686_ (.A1(_0367_),
    .A2(_0377_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2687_ (.A1(_0215_),
    .A2(_0214_),
    .A3(_0269_),
    .A4(_0341_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2688_ (.A1(_0193_),
    .A2(_0379_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2689_ (.I(_0059_),
    .Z(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2690_ (.I(_0182_),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2691_ (.A1(_0046_),
    .A2(_0033_),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2692_ (.A1(_0105_),
    .A2(_0221_),
    .Z(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2693_ (.A1(_0324_),
    .A2(_1416_),
    .B1(_0384_),
    .B2(_0383_),
    .C(_0385_),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2694_ (.A1(_0383_),
    .A2(_0384_),
    .A3(_0385_),
    .B(_0386_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2695_ (.A1(_0381_),
    .A2(_0387_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2696_ (.A1(_0121_),
    .A2(_0336_),
    .B(_0388_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2697_ (.A1(_0380_),
    .A2(_0389_),
    .Z(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2698_ (.I(_0052_),
    .Z(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2699_ (.A1(_0324_),
    .A2(_1415_),
    .A3(_0033_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2700_ (.A1(_0391_),
    .A2(_0136_),
    .B(_0392_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2701_ (.A1(_0100_),
    .A2(_0292_),
    .A3(_0293_),
    .A4(_0384_),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2702_ (.A1(_0324_),
    .A2(_0323_),
    .A3(_0181_),
    .B(_0381_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2703_ (.A1(_1315_),
    .A2(_1340_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2704_ (.A1(_0288_),
    .A2(_0397_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2705_ (.A1(_0394_),
    .A2(_0395_),
    .A3(_0396_),
    .B1(_0398_),
    .B2(_0381_),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2706_ (.A1(_0162_),
    .A2(_0399_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2707_ (.A1(_0279_),
    .A2(_0400_),
    .Z(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2708_ (.A1(_0115_),
    .A2(_0390_),
    .A3(_0401_),
    .Z(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2709_ (.A1(_0115_),
    .A2(_0390_),
    .B(_0401_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2710_ (.A1(_0114_),
    .A2(_0402_),
    .A3(_0403_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2711_ (.A1(_0378_),
    .A2(_0405_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _2712_ (.A1(_0366_),
    .A2(_0406_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2713_ (.A1(_0173_),
    .A2(_0231_),
    .B(_0313_),
    .C(_0356_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2714_ (.A1(_0319_),
    .A2(_0355_),
    .Z(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2715_ (.A1(_0319_),
    .A2(_0355_),
    .Z(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2716_ (.A1(_0360_),
    .A2(_0409_),
    .B(_0410_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2717_ (.A1(_0310_),
    .A2(_0408_),
    .B(_0411_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2718_ (.A1(_0407_),
    .A2(_0412_),
    .Z(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2719_ (.I(_0413_),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2720_ (.A1(_0378_),
    .A2(_0405_),
    .B(_0402_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2721_ (.I(_0166_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2722_ (.A1(_0369_),
    .A2(_1361_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _2723_ (.A1(_0293_),
    .A2(_1375_),
    .B(_0185_),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2724_ (.A1(_0054_),
    .A2(_0369_),
    .B(_0417_),
    .C(_0418_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2725_ (.A1(_0284_),
    .A2(_0294_),
    .A3(_0259_),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2726_ (.A1(_0368_),
    .A2(_0419_),
    .B(_0420_),
    .C(_0283_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2727_ (.A1(_0380_),
    .A2(_0421_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2728_ (.A1(_0062_),
    .A2(_0343_),
    .B(_0342_),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2729_ (.A1(_0197_),
    .A2(_0418_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2730_ (.A1(_0262_),
    .A2(_0323_),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2731_ (.A1(_0285_),
    .A2(_0044_),
    .B(_0426_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2732_ (.A1(_0131_),
    .A2(_1327_),
    .B(_0174_),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2733_ (.A1(_0132_),
    .A2(_0428_),
    .B(_0282_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _2734_ (.A1(_0208_),
    .A2(_0424_),
    .B1(_0427_),
    .B2(_0184_),
    .C(_0429_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2735_ (.A1(_1428_),
    .A2(_0430_),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2736_ (.A1(_0423_),
    .A2(_0430_),
    .B(_0431_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2737_ (.A1(_0162_),
    .A2(_0432_),
    .Z(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2738_ (.A1(_0416_),
    .A2(_0422_),
    .B(_0433_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2739_ (.A1(_0416_),
    .A2(_0433_),
    .A3(_0422_),
    .Z(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2740_ (.A1(_0232_),
    .A2(_0434_),
    .A3(_0435_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2741_ (.I(_0367_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2742_ (.A1(_0375_),
    .A2(_1422_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2743_ (.I(_1372_),
    .Z(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2744_ (.A1(_0391_),
    .A2(_0203_),
    .A3(_0204_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2745_ (.A1(_0440_),
    .A2(_1416_),
    .A3(_0441_),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2746_ (.A1(_0133_),
    .A2(_0442_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2747_ (.A1(_0289_),
    .A2(_0439_),
    .B1(_0443_),
    .B2(_0375_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2748_ (.A1(_0438_),
    .A2(_0444_),
    .Z(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2749_ (.A1(_0437_),
    .A2(_0445_),
    .Z(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _2750_ (.A1(_0415_),
    .A2(_0446_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2751_ (.A1(_0366_),
    .A2(_0406_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2752_ (.A1(_0407_),
    .A2(_0412_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2753_ (.A1(_0449_),
    .A2(_0450_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2754_ (.A1(_0448_),
    .A2(_0451_),
    .Z(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2755_ (.I(_0452_),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2756_ (.A1(_0437_),
    .A2(_0445_),
    .B(_0435_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2757_ (.A1(_0284_),
    .A2(_0078_),
    .A3(_0197_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2758_ (.A1(_1372_),
    .A2(_1293_),
    .A3(_1440_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2759_ (.A1(_0283_),
    .A2(_0454_),
    .A3(_0455_),
    .B1(_1432_),
    .B2(_0426_),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2760_ (.A1(_0368_),
    .A2(_1285_),
    .A3(_0073_),
    .B(_0456_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2761_ (.I0(_0063_),
    .I1(_0423_),
    .S(_0458_),
    .Z(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2762_ (.A1(_0350_),
    .A2(_0432_),
    .B(_1390_),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2763_ (.A1(_0350_),
    .A2(_0459_),
    .B(_0460_),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2764_ (.I(_0368_),
    .Z(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2765_ (.A1(_0273_),
    .A2(_0418_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2766_ (.A1(_0462_),
    .A2(_0463_),
    .ZN(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2767_ (.A1(_1364_),
    .A2(_0323_),
    .B(_0321_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2768_ (.A1(_0381_),
    .A2(_0464_),
    .A3(_0465_),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2769_ (.A1(_0291_),
    .A2(_0379_),
    .B(_0193_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2770_ (.A1(_0466_),
    .A2(_0467_),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2771_ (.A1(_0267_),
    .A2(_0466_),
    .B(_0469_),
    .C(_0416_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2772_ (.A1(_0461_),
    .A2(_0470_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2773_ (.A1(_0328_),
    .A2(_0330_),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2774_ (.A1(_0097_),
    .A2(_0218_),
    .B1(_0248_),
    .B2(_0391_),
    .C(_0462_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2775_ (.A1(_0472_),
    .A2(_0473_),
    .B(_0233_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2776_ (.I0(_0233_),
    .I1(_0474_),
    .S(_0611_),
    .Z(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2777_ (.A1(_0471_),
    .A2(_0475_),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2778_ (.A1(_0453_),
    .A2(_0476_),
    .Z(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2779_ (.A1(_0415_),
    .A2(_0446_),
    .B(_0449_),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2780_ (.A1(_0415_),
    .A2(_0446_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2781_ (.A1(_0407_),
    .A2(_0412_),
    .A3(_0448_),
    .B1(_0478_),
    .B2(_0480_),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2782_ (.A1(_0477_),
    .A2(_0481_),
    .Z(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2783_ (.I(_0482_),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2784_ (.A1(_0461_),
    .A2(_0470_),
    .Z(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2785_ (.A1(_0471_),
    .A2(_0475_),
    .B(_0483_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2786_ (.I(_0484_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2787_ (.I(_0374_),
    .Z(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2788_ (.A1(_0486_),
    .A2(_0080_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2789_ (.A1(_0146_),
    .A2(_0222_),
    .A3(_0487_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2790_ (.I0(_0611_),
    .I1(_0438_),
    .S(_0488_),
    .Z(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2791_ (.I(_0369_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2792_ (.A1(_0491_),
    .A2(_0176_),
    .ZN(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2793_ (.A1(_0492_),
    .A2(_1440_),
    .B(_1329_),
    .C(_1437_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2794_ (.A1(_0096_),
    .A2(_0273_),
    .B1(_0473_),
    .B2(_0375_),
    .C(_0493_),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2795_ (.A1(_0063_),
    .A2(_0494_),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2796_ (.A1(_0280_),
    .A2(_0494_),
    .B(_0495_),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2797_ (.A1(_0350_),
    .A2(_0496_),
    .B(_0460_),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2798_ (.A1(_0080_),
    .A2(_0383_),
    .B(_0440_),
    .ZN(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2799_ (.A1(_0440_),
    .A2(_0418_),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2800_ (.A1(_0374_),
    .A2(_0499_),
    .ZN(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2801_ (.A1(_0498_),
    .A2(_0501_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2802_ (.A1(_0380_),
    .A2(_0502_),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2803_ (.A1(_0267_),
    .A2(_0502_),
    .B(_0503_),
    .C(_0234_),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2804_ (.A1(_0497_),
    .A2(_0504_),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2805_ (.A1(_0497_),
    .A2(_0504_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2806_ (.A1(_0505_),
    .A2(_0506_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2807_ (.A1(_0490_),
    .A2(_0507_),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2808_ (.A1(_0453_),
    .A2(_0476_),
    .Z(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2809_ (.A1(_0477_),
    .A2(_0481_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2810_ (.A1(_0509_),
    .A2(_0510_),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2811_ (.A1(_0485_),
    .A2(_0508_),
    .A3(_0512_),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2812_ (.I(_0513_),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2813_ (.A1(_0285_),
    .A2(_1407_),
    .B(_0325_),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2814_ (.A1(_0109_),
    .A2(_0337_),
    .B1(_0514_),
    .B2(_0374_),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2815_ (.A1(_0148_),
    .A2(_0279_),
    .Z(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2816_ (.A1(_0515_),
    .A2(_0516_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2817_ (.A1(_0025_),
    .A2(_0517_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2818_ (.A1(_0462_),
    .A2(_1429_),
    .B(_0501_),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2819_ (.A1(_0380_),
    .A2(_0519_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _2820_ (.A1(_0267_),
    .A2(_0519_),
    .B(_0520_),
    .C(_0416_),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2821_ (.A1(_0518_),
    .A2(_0522_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2822_ (.A1(_0610_),
    .A2(_0222_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2823_ (.A1(_0222_),
    .A2(_0367_),
    .B(_0524_),
    .C(_0146_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2824_ (.I(_0525_),
    .Z(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2825_ (.A1(_0523_),
    .A2(_0526_),
    .Z(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2826_ (.A1(_0490_),
    .A2(_0507_),
    .B(_0505_),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2827_ (.A1(_0527_),
    .A2(_0528_),
    .Z(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2828_ (.A1(_0485_),
    .A2(_0508_),
    .Z(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2829_ (.A1(_0485_),
    .A2(_0508_),
    .B(_0509_),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2830_ (.A1(_0477_),
    .A2(_0481_),
    .B(_0531_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2831_ (.A1(_0530_),
    .A2(_0533_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2832_ (.A1(_0529_),
    .A2(_0534_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2833_ (.I(_0535_),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2834_ (.A1(_0518_),
    .A2(_0522_),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2835_ (.A1(_0523_),
    .A2(_0526_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2836_ (.A1(_0391_),
    .A2(_1407_),
    .B(_0109_),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2837_ (.A1(_0370_),
    .A2(_0462_),
    .B(_0486_),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2838_ (.A1(_0538_),
    .A2(_0539_),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2839_ (.A1(_0280_),
    .A2(_0540_),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2840_ (.A1(_0063_),
    .A2(_0540_),
    .B(_0541_),
    .ZN(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2841_ (.A1(_0159_),
    .A2(_0543_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2842_ (.A1(_0460_),
    .A2(_0544_),
    .Z(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2843_ (.A1(_0522_),
    .A2(_0525_),
    .A3(_0545_),
    .Z(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2844_ (.A1(_0536_),
    .A2(_0537_),
    .B(_0546_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2845_ (.A1(_0536_),
    .A2(_0537_),
    .A3(_0546_),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2846_ (.A1(_0547_),
    .A2(_0548_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2847_ (.I(_0529_),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2848_ (.A1(_0527_),
    .A2(_0528_),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2849_ (.A1(_0530_),
    .A2(_0550_),
    .A3(_0533_),
    .B(_0551_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2850_ (.A1(_0549_),
    .A2(_0552_),
    .Z(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2851_ (.I(_0554_),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2852_ (.A1(_0526_),
    .A2(_0545_),
    .ZN(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2853_ (.A1(_0526_),
    .A2(_0545_),
    .B(_0522_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2854_ (.A1(_0555_),
    .A2(_0556_),
    .ZN(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2855_ (.A1(_0529_),
    .A2(_0549_),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2856_ (.A1(_0530_),
    .A2(_0533_),
    .A3(_0558_),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2857_ (.A1(_0536_),
    .A2(_0537_),
    .A3(_0546_),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2858_ (.A1(_0551_),
    .A2(_0560_),
    .B(_0547_),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _2859_ (.A1(_0557_),
    .A2(_0559_),
    .A3(_0561_),
    .B1(_0516_),
    .B2(_0232_),
    .ZN(net7));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2860_ (.A1(_1396_),
    .A2(_0089_),
    .Z(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2861_ (.I(_0563_),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2862_ (.A1(\bit2symb.regi ),
    .A2(_0265_),
    .ZN(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2863_ (.A1(_0611_),
    .A2(net42),
    .B(_0564_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2864_ (.I0(\Reg_Delay_Q.In ),
    .I1(net1),
    .S(_0265_),
    .Z(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2865_ (.I(_0565_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2866_ (.A1(_0383_),
    .A2(_0439_),
    .ZN(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2867_ (.I(_0566_),
    .Z(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2868_ (.A1(\Reg_Delay_Q.In ),
    .A2(_0567_),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2869_ (.A1(_0619_),
    .A2(_0567_),
    .B(_0568_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2870_ (.I(net2),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2871_ (.A1(_1399_),
    .A2(_0570_),
    .Z(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2872_ (.I(_0571_),
    .Z(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2873_ (.I(_0570_),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2874_ (.A1(_0570_),
    .A2(_0176_),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2875_ (.A1(_1277_),
    .A2(_0572_),
    .B1(net44),
    .B2(_0573_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2876_ (.A1(net2),
    .A2(_1361_),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2877_ (.A1(_0491_),
    .A2(_0574_),
    .Z(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2878_ (.I(_0575_),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2879_ (.A1(_0491_),
    .A2(_0574_),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2880_ (.A1(_0370_),
    .A2(_0576_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2881_ (.I(_0578_),
    .Z(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2882_ (.A1(_0370_),
    .A2(_0576_),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2883_ (.A1(_0203_),
    .A2(_1422_),
    .B(_0609_),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2884_ (.A1(_0440_),
    .A2(_0579_),
    .B1(_0580_),
    .B2(_0572_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2885_ (.A1(_0491_),
    .A2(_1422_),
    .A3(_0574_),
    .ZN(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2886_ (.I(net2),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2887_ (.I(_0582_),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2888_ (.A1(_0583_),
    .A2(_0133_),
    .B1(_0581_),
    .B2(_0486_),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2889_ (.A1(_0486_),
    .A2(_0581_),
    .B(_0584_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2890_ (.A1(_0582_),
    .A2(_0567_),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2891_ (.I(_0586_),
    .Z(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2892_ (.A1(_0844_),
    .A2(_0583_),
    .ZN(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2893_ (.A1(_0844_),
    .A2(_0587_),
    .B(_0588_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2894_ (.A1(_0647_),
    .A2(_0572_),
    .B1(_0663_),
    .B2(_0587_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2895_ (.A1(_0763_),
    .A2(_0755_),
    .A3(_0587_),
    .B1(_0572_),
    .B2(_1075_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2896_ (.A1(_1038_),
    .A2(_0774_),
    .A3(_0586_),
    .B1(_0570_),
    .B2(_0809_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2897_ (.A1(_0582_),
    .A2(_0775_),
    .A3(_0566_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2898_ (.A1(_0582_),
    .A2(_0589_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2899_ (.A1(_1227_),
    .A2(_0590_),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2900_ (.A1(_0889_),
    .A2(_0653_),
    .A3(_0589_),
    .B(_0591_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2901_ (.A1(_1202_),
    .A2(_0590_),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2902_ (.A1(_1202_),
    .A2(_0775_),
    .A3(_0587_),
    .B(_0593_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2903_ (.A1(_1122_),
    .A2(\p_shaping_Q.counter[0] ),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2904_ (.A1(_0022_),
    .A2(_0594_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2905_ (.A1(_0609_),
    .A2(_0567_),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2906_ (.I0(\bit2symb.regi ),
    .I1(net1),
    .S(_0595_),
    .Z(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2907_ (.I(_0596_),
    .Z(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2908_ (.A1(_0234_),
    .A2(\p_shaping_I.counter[0] ),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2909_ (.A1(_0025_),
    .A2(_0597_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2910_ (.D(_0006_),
    .RN(net63),
    .CLK(clknet_1_1__leaf_CLK),
    .Q(\p_shaping_I.bit_in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2911_ (.D(_0007_),
    .RN(net60),
    .CLK(clknet_1_1__leaf_CLK),
    .Q(\Reg_Delay_Q.In ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2912_ (.D(_0008_),
    .RN(net63),
    .CLK(clknet_1_1__leaf_CLK),
    .Q(\Reg_Delay_Q.Out ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2913_ (.D(_0009_),
    .RN(net56),
    .CLK(clknet_1_0__leaf_CLK),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2914_ (.D(_0010_),
    .RN(net57),
    .CLK(clknet_1_0__leaf_CLK),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2915_ (.D(_0011_),
    .RN(net56),
    .CLK(clknet_1_0__leaf_CLK),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2916_ (.D(_0012_),
    .RN(net58),
    .CLK(clknet_1_0__leaf_CLK),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _2917_ (.D(_0013_),
    .RN(net59),
    .CLK(clknet_1_1__leaf_CLK),
    .Q(net34));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _2918_ (.D(_0014_),
    .RN(net60),
    .CLK(clknet_1_1__leaf_CLK),
    .Q(net35));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2919_ (.D(_0015_),
    .RN(net57),
    .CLK(clknet_1_0__leaf_CLK),
    .Q(net36));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2920_ (.D(_0016_),
    .RN(net56),
    .CLK(clknet_1_0__leaf_CLK),
    .Q(net37));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2921_ (.D(_0017_),
    .RN(net56),
    .CLK(clknet_1_0__leaf_CLK),
    .Q(net38));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2922_ (.D(_0018_),
    .RN(net58),
    .CLK(clknet_1_0__leaf_CLK),
    .Q(net39));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _2923_ (.D(_0019_),
    .RN(net58),
    .CLK(clknet_1_0__leaf_CLK),
    .Q(net40));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2924_ (.D(_0020_),
    .RN(net60),
    .CLK(clknet_1_1__leaf_CLK),
    .Q(net41));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2925_ (.D(_0021_),
    .RN(net61),
    .CLK(net48),
    .Q(\p_shaping_Q.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2926_ (.D(_0022_),
    .RN(net62),
    .CLK(net48),
    .Q(\p_shaping_Q.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__latrnq_1 _2927_ (.D(_0000_),
    .Q(\p_shaping_I.ctl_1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2928_ (.D(\p_shaping_I.bit_in ),
    .RN(net61),
    .CLK(net42),
    .Q(\p_shaping_I.bit_in_1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2929_ (.D(\p_shaping_I.bit_in_1 ),
    .RN(net65),
    .CLK(net42),
    .Q(\p_shaping_I.bit_in_2 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2930_ (.D(_0023_),
    .RN(net60),
    .CLK(clknet_1_1__leaf_CLK),
    .Q(\bit2symb.regi ));
 gf180mcu_fd_sc_mcu7t5v0__latrnq_1 _2931_ (.D(_0002_),
    .Q(\p_shaping_Q.ctl_1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2932_ (.D(\Reg_Delay_Q.Out ),
    .RN(net63),
    .CLK(net47),
    .Q(\p_shaping_Q.bit_in_1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2933_ (.D(\p_shaping_Q.bit_in_1 ),
    .RN(net62),
    .CLK(net48),
    .Q(\p_shaping_Q.bit_in_2 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2934_ (.D(_0024_),
    .RN(net61),
    .CLK(net43),
    .Q(\p_shaping_I.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2935_ (.D(_0025_),
    .RN(net61),
    .CLK(net43),
    .Q(\p_shaping_I.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_CLK (.I(CLK),
    .Z(clknet_0_CLK));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_0__f_CLK (.I(clknet_0_CLK),
    .Z(clknet_1_0__leaf_CLK));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_1__f_CLK (.I(clknet_0_CLK),
    .Z(clknet_1_1__leaf_CLK));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout42 (.I(net44),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout43 (.I(net44),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout44 (.I(_0004_),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout47 (.I(_0005_),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout48 (.I(_0005_),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout49 (.I(net41),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout50 (.I(net39),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout51 (.I(net37),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout52 (.I(net36),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout53 (.I(net33),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout54 (.I(net31),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout55 (.I(net30),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout56 (.I(net57),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout57 (.I(net58),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout58 (.I(net59),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout59 (.I(net66),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout60 (.I(net65),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout61 (.I(net64),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout62 (.I(net64),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout63 (.I(net65),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout64 (.I(net65),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout65 (.I(net66),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout66 (.I(net3),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1 (.I(BitIn),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(EN),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(RST),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output10 (.I(net10),
    .Z(I[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output11 (.I(net11),
    .Z(I[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output12 (.I(net12),
    .Z(I[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output13 (.I(net13),
    .Z(I[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output14 (.I(net14),
    .Z(I[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output15 (.I(net15),
    .Z(I[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output16 (.I(net16),
    .Z(I[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output17 (.I(net17),
    .Z(Q[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output18 (.I(net18),
    .Z(Q[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output19 (.I(net19),
    .Z(Q[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output20 (.I(net20),
    .Z(Q[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output21 (.I(net21),
    .Z(Q[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output22 (.I(net22),
    .Z(Q[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output23 (.I(net23),
    .Z(Q[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output24 (.I(net24),
    .Z(Q[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output25 (.I(net25),
    .Z(Q[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output26 (.I(net26),
    .Z(Q[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output27 (.I(net27),
    .Z(Q[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output28 (.I(net28),
    .Z(Q[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output29 (.I(net29),
    .Z(Q[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output30 (.I(net55),
    .Z(addI[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output31 (.I(net54),
    .Z(addI[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output32 (.I(net32),
    .Z(addI[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output33 (.I(net53),
    .Z(addI[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output34 (.I(net34),
    .Z(addI[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output35 (.I(net35),
    .Z(addI[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output36 (.I(net52),
    .Z(addQ[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output37 (.I(net51),
    .Z(addQ[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output38 (.I(net38),
    .Z(addQ[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output39 (.I(net39),
    .Z(addQ[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output4 (.I(net4),
    .Z(I[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output40 (.I(net40),
    .Z(addQ[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output41 (.I(net41),
    .Z(addQ[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output5 (.I(net5),
    .Z(I[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output6 (.I(net6),
    .Z(I[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output7 (.I(net7),
    .Z(I[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output8 (.I(net8),
    .Z(I[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output9 (.I(net9),
    .Z(I[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wire45 (.I(_0299_),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wire46 (.I(_1100_),
    .Z(net46));
 assign io_oeb[0] = net98;
 assign io_oeb[10] = net70;
 assign io_oeb[11] = net71;
 assign io_oeb[12] = net72;
 assign io_oeb[13] = net73;
 assign io_oeb[14] = net74;
 assign io_oeb[15] = net75;
 assign io_oeb[16] = net76;
 assign io_oeb[17] = net77;
 assign io_oeb[18] = net78;
 assign io_oeb[19] = net79;
 assign io_oeb[1] = net99;
 assign io_oeb[20] = net80;
 assign io_oeb[21] = net81;
 assign io_oeb[22] = net82;
 assign io_oeb[23] = net83;
 assign io_oeb[24] = net84;
 assign io_oeb[25] = net85;
 assign io_oeb[26] = net86;
 assign io_oeb[27] = net87;
 assign io_oeb[28] = net88;
 assign io_oeb[29] = net89;
 assign io_oeb[2] = net100;
 assign io_oeb[30] = net90;
 assign io_oeb[31] = net91;
 assign io_oeb[32] = net92;
 assign io_oeb[33] = net93;
 assign io_oeb[34] = net94;
 assign io_oeb[35] = net95;
 assign io_oeb[36] = net96;
 assign io_oeb[37] = net97;
 assign io_oeb[3] = net101;
 assign io_oeb[4] = net102;
 assign io_oeb[5] = net103;
 assign io_oeb[6] = net104;
 assign io_oeb[7] = net67;
 assign io_oeb[8] = net68;
 assign io_oeb[9] = net69;
endmodule

