* NGSPICE file created from OQPSK_PS_RCOSINE2.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 D RN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__latrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__latrnq_1 D E RN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_1 A1 A2 A3 B1 B2 B3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_4 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_2 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VNW VPW VSS
.ends

.subckt OQPSK_PS_RCOSINE2 BitIn CLK EN I[0] I[10] I[11] I[12] I[1] I[2] I[3] I[4]
+ I[5] I[6] I[7] I[8] I[9] Q[0] Q[10] Q[11] Q[12] Q[1] Q[2] Q[3] Q[4] Q[5] Q[6] Q[7]
+ Q[8] Q[9] RST addI[0] addI[1] addI[2] addI[3] addI[4] addI[5] addQ[0] addQ[1] addQ[2]
+ addQ[3] addQ[4] addQ[5] io_oeb[0] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[2] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3]
+ io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] vdd vss io_oeb[29] io_oeb[28]
+ io_oeb[27] io_oeb[26] io_oeb[25] io_oeb[13] io_oeb[24] io_oeb[23] io_oeb[12] io_oeb[33]
+ io_oeb[22] io_oeb[11] io_oeb[21] io_oeb[10] io_oeb[32] io_oeb[20] io_oeb[31] io_oeb[30]
X_2106_ _1104_ _1176_ _1177_ _0670_ _1178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_2037_ _0730_ _1108_ _1110_ _0672_ _1111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_49_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1606_ net49 _0684_ _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_54_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2724_ _0054_ _0369_ _0417_ _0418_ _0419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_14_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2655_ _0333_ _0341_ _1323_ _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2164__A2 _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1537_ Reg_Delay_Q.Out _0619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_1468_ net34 _0124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_1_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2586_ _1400_ _0107_ _0181_ _0272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__1675__A1 _0752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_56_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_5_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2440_ _1391_ _0114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_11_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2371_ _1372_ _0032_ _0037_ _0038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__2449__A3 _1366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2909__A1 _0025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2137__A2 _0663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2638_ _0282_ _1429_ _0326_ _0327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2385__A2 _1314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2707_ _0279_ _0400_ _0401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2569_ _0188_ _0111_ _0187_ _0253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_65_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1648__A1 _0700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1820__A1 _0887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2300__A2 _1375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1940_ _0907_ _0956_ _0957_ _1016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1871_ _0542_ _0892_ _0948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_43_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2423_ _1322_ _1411_ _0094_ _0095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2367__A2 _1337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2285_ _1353_ _1286_ _1360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2354_ _1309_ _1351_ _1434_ _1435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2294__A1 _1367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1487__I _0318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_13_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1950__I _0852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2070_ _0618_ _1141_ _1094_ _1143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XPHY_EDGE_ROW_28_Left_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1854_ _0748_ _0911_ _0746_ _0704_ _0931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_1785_ p_shaping_Q.bit_in_1 _0863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1923_ _0854_ _0890_ _0772_ _0812_ _0999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__2588__A2 _0273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2760__A2 _1285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2406_ _1335_ _1286_ _1295_ _0076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_2199_ _1242_ _1259_ _1235_ _1267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2268_ _0211_ _0124_ _1341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_2337_ _1298_ _1326_ _1300_ _1416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_43_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2503__A2 _1375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1570_ _0648_ _0649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2742__A2 _1422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2122_ _1189_ _1193_ _0619_ _1194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2053_ _0808_ _1126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_16_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1906_ _0839_ _0768_ _0981_ _0923_ _0982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_1768_ _0656_ _0843_ _0845_ _0846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1837_ _0742_ _0659_ _0914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2886_ net2 _0582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2430__A1 _0101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1699_ _0692_ _0643_ _0678_ _0777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_0_67_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput20 net20 Q[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput31 net54 addI[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput7 net7 I[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__2724__A2 _0369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1714__B _0791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1622_ p_shaping_Q.counter\[1\] _0701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2740_ _0232_ _0434_ _0435_ _0437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_2671_ _0360_ _0362_ _0363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1484_ _0286_ _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1553_ net51 _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout49_I net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2105_ _1104_ _0998_ _1177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_2036_ _1109_ _1103_ _0942_ _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_37_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2921__CLK clknet_1_0__leaf_CLK vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2869_ _0619_ _0567_ _0568_ _0008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_4_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2706__A2 _0399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_15_Left_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2642__A1 _0328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_59_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2723_ _0293_ _1375_ _0185_ _0418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_1536_ _0617_ _0618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1605_ _0318_ _0675_ _0340_ _0414_ _0684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2585_ _0234_ _0266_ _0270_ _0271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2654_ _0342_ _0343_ _0344_ _0149_ _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_1467_ _0102_ _0113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__1978__A3 _1051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2019_ _1083_ _1092_ _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_9_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_0_Left_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1666__A2 _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2863__A1 _0611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2370_ _1402_ _1417_ _1307_ _0037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_59_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2706_ _0162_ _0399_ _0400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2733__B _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1519_ net49 _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2637_ _0323_ _0221_ _0325_ _0326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2568_ _0096_ _0245_ _0246_ _0247_ _0251_ _0252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2499_ _0175_ _0176_ _0064_ _1374_ _0130_ _0177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_36_Left_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_45_Left_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2300__A3 _1369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1870_ _0598_ _0718_ _0947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_EDGE_ROW_54_Left_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_63_Left_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1575__B2 _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2422_ p_shaping_I.bit_in _0094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2353_ _1306_ _1362_ _1433_ _1434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_19_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2284_ _1358_ _1359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1999_ _1031_ _1072_ _1073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_30_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2689__I _0059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2530__A3 _0127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_3_Left_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1922_ _0864_ _0997_ _0616_ _0998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_56_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1784_ _0669_ _0862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1853_ _0926_ _0929_ _0930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_44_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2405_ _1404_ _0048_ _0049_ _0075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__2760__A3 _0073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2336_ _1353_ _1343_ _1441_ _1415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_67_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2198_ _1242_ _1259_ _1266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2267_ _1305_ _1289_ _1336_ _1340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_62_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2019__A2 _1092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2121_ _1072_ _1192_ _1189_ _1193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2052_ _1079_ _1125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1905_ _0828_ _0858_ _0846_ _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2885_ _0491_ _1422_ _0574_ _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__2430__A2 _1340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1698_ _0703_ _0748_ _0773_ _0674_ _0775_ _0776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_1767_ _0844_ _0817_ _0748_ _0845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1836_ _0740_ _0649_ _0637_ _0913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_25_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2319_ _1392_ _1395_ _1396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_67_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput21 net21 Q[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput32 net32 addI[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__2327__I3 _1403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput8 net8 I[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput10 net10 I[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XPHY_EDGE_ROW_59_Right_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_46_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2561__B _0221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1621_ _0674_ _0686_ _0690_ _0696_ _0698_ _0699_ _0700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_1552_ _0630_ _0631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2670_ _0310_ _0314_ _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2104_ _1057_ _1174_ _1175_ _1176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1483_ net52 _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input3_I RST vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2035_ _0997_ _1059_ _0863_ _1109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__2100__B2 _0927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_37_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2190__C _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2868_ Reg_Delay_Q.In _0567_ _0568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1819_ _0891_ _0892_ _0894_ _0896_ _0639_ _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__1914__A1 _0308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2799_ _0440_ _0418_ _0499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2330__A1 _1296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2722_ _0369_ _1361_ _0417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1535_ _0616_ _0617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1604_ _0681_ _0682_ _0635_ _0683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_0_1_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2584_ _0267_ _0268_ _0269_ _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2653_ _1428_ _0278_ _0344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_38_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1466_ _1258_ _1354_ _0102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_49_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2018_ _0771_ _1089_ _1091_ _0500_ _1092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_45_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2823__C _0146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2551__A1 _0234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_19_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2636_ _0185_ _0293_ _0324_ _0325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2705_ _0394_ _0395_ _0396_ _0398_ _0381_ _0399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_6_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1518_ _0599_ _0601_ _0602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_49_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2498_ _1313_ _0176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_2_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2567_ _0185_ _0248_ _0249_ _0250_ _0121_ _0251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1449_ _1321_ _1332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2533__A1 _0199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_43_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2421_ _0092_ _0088_ _0087_ _0093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2283_ _1289_ _1358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2352_ _1295_ _1433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_19_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1998_ _0980_ _0982_ _1030_ _1072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_30_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2619_ _0304_ _0306_ _0232_ _0307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_15_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2818__A2 _1429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2294__A3 _1369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1784__I _0669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1921_ _0873_ _0877_ _0945_ _0950_ _0997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_56_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1852_ _0927_ _0928_ _0929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1796__A2 _0777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1783_ _0841_ _0860_ _0861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_52_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2745__A1 _0440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2335_ p_shaping_I.bit_in_2 _1330_ _1334_ _1342_ _1414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_2266_ _1331_ _1338_ _1339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2404_ _0071_ _0073_ _0034_ _0074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2197_ _1265_ net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2120_ _1078_ _1190_ _1191_ _1192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_21_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2051_ _0960_ _1082_ _1107_ _1123_ _1124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_16_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1835_ _0817_ _0911_ _0912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1904_ _0973_ _0979_ _0980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2884_ _0440_ _0579_ _0580_ _0572_ _0013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_32_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1766_ _0308_ _0844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1697_ _0673_ _0774_ _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__2313__I _1390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2318_ _1322_ _1393_ _1395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2249_ _1279_ _1304_ _1319_ _0146_ _1320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__1457__A1 net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2223__I _0091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput22 net22 Q[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__1932__A2 _1001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput33 net53 addI[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_31_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput9 net9 I[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput11 net11 I[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_58_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1620_ _0685_ _0699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1551_ _0626_ _0629_ _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_41_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1482_ _0265_ _0004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2289__B _1363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2103_ _0863_ _1174_ _1175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_37_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2034_ _1083_ _1092_ _1108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_49_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1818_ _0740_ _0707_ _0697_ _0797_ _0895_ _0896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__1611__A1 _0687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2867_ _0566_ _0567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2798_ _0080_ _0383_ _0440_ _0498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1749_ _0650_ _0826_ _0732_ _0827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1831__B _0752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2875__B1 net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1669__A1 _0647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2837__B _0486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1841__B2 _0852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2721_ _0166_ _0416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2652_ _0278_ _0343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_1534_ p_shaping_Q.bit_in_1 _0616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1603_ _0340_ _0682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1465_ net53 _0091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_22_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2583_ _0258_ _0261_ _0263_ _0269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_2017_ _1090_ _0754_ _1091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_65_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2919_ _0015_ net57 clknet_1_0__leaf_CLK net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_9_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2501__I _1416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output35_I net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2303__A2 _1366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2067__A1 _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2635_ _1406_ _0324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2704_ _0288_ _0397_ _0398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1517_ _0468_ _0600_ _0601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1448_ net55 _1321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2566_ _0100_ _1359_ _0250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2497_ _1285_ _0175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1805__A1 _0705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2297__A1 _1357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2420_ _1413_ _0092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_3_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2351_ _1278_ _1431_ _1432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_2282_ _1355_ _1294_ _1356_ _1357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_59_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1997_ _1033_ _1065_ _1063_ _1071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_51_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2460__A1 _1417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2618_ _0159_ _0301_ _0305_ _0306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_15_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2549_ _1390_ _0232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_38_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2451__A1 _0108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1920_ _0985_ _0986_ _0994_ _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_56_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1851_ _0635_ _0716_ _0928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_37_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1782_ _0846_ _0859_ _0860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2745__A2 _1416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2403_ _1355_ _0072_ _1290_ _0073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_12_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2196_ _1263_ _1264_ _1265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2334_ _1411_ _1412_ _1413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2265_ _1335_ _1282_ _1365_ _1338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_47_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2736__A2 _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2649__C _1406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2050_ _1122_ _1093_ _1106_ _1123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2575__B _0136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1765_ _0743_ _0710_ _0842_ _0843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1834_ _0910_ _0911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1903_ _0974_ _0977_ _0978_ _0948_ _0828_ _0979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_44_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2883_ _0203_ _1422_ _0609_ _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_32_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1696_ _0425_ _0652_ _0774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_57_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2179_ _1245_ _1247_ _1248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_2317_ _1394_ net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2248_ _1309_ _1315_ _1318_ _1319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput23 net23 Q[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput34 net34 addI[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput12 net12 I[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__2893__A1 _0844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1550_ _0628_ _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1481_ _0254_ _0265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2102_ _1074_ _0646_ _0933_ _1169_ _1173_ _1174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_2033_ _0925_ _1093_ _1106_ _1107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_37_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2884__A1 _0440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2935_ _0025_ net61 net43 p_shaping_I.counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_9_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1817_ _0762_ _0711_ _0895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1748_ _0382_ _0781_ _0351_ _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_25_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2866_ _0383_ _0439_ _0566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2797_ _0350_ _0496_ _0460_ _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1679_ _0755_ _0756_ _0757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1678__A2 _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2875__A1 _1277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1669__A2 _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2866__A1 _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1602_ _0675_ _0681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2651_ _0155_ _0225_ _0607_ _0342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_1_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2720_ _0378_ _0405_ _0402_ _0415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2582_ _0210_ _0212_ _0268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1464_ _1441_ _0069_ _1288_ _0080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1533_ _0608_ _0609_ _0615_ _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_65_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2016_ _0812_ _1090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_19_Left_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2918_ _0014_ net60 clknet_1_1__leaf_CLK net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2849_ _0530_ _0550_ _0533_ _0551_ _0552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__1520__A1 _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2567__C _0121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1516_ _0361_ _0600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2703_ _1315_ _1340_ _0397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_2_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2565_ _0055_ _1361_ _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2634_ _0064_ _0323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_65_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2496_ _0130_ _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1447_ _1299_ _1310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__1805__A2 _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1741__A1 _0818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2297__A2 _1364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_32_Left_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2350_ _1317_ _1429_ _1431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2281_ _1307_ _1356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_19_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1996_ _1070_ net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1723__A1 _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2617_ _0149_ _0279_ _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2548_ _0191_ _0230_ _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_2479_ _0155_ _0156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_65_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2451__A2 _1415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1781_ _0822_ _0858_ _0859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_56_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1850_ _0479_ _0759_ _0927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1705__A1 _0742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2333_ p_shaping_I.bit_in _1322_ _1412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2402_ _1332_ _0072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_46_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2195_ _1222_ _1248_ _1251_ _1245_ _1247_ _1264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_27_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2264_ _1335_ _1336_ _1337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_47_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1979_ _1049_ _1052_ _0733_ _1053_ _1054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_43_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_7_Left_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2112__A1 _1001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2575__C _0051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1902_ _0971_ _0975_ _0819_ _0978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_32_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1764_ _0793_ _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1833_ _0633_ _0297_ _0678_ _0910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_40_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2882_ _0370_ _0576_ _0579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_32_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1695_ _0720_ _0772_ _0636_ _0630_ _0773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_2316_ _1322_ _1393_ _1394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_12_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2178_ _1207_ _1219_ _1246_ _1247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2247_ _1316_ _1317_ _1318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__1917__A1 _0887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput24 net24 Q[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_31_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput35 net35 addI[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput13 net13 I[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_16_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2645__A2 _0181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1480_ _0243_ _0254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2586__B _0181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2101_ _0928_ _1170_ _1172_ _0808_ _1029_ _1173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_2032_ _1094_ _1103_ _1105_ _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_37_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2914__CLK clknet_1_0__leaf_CLK vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2865_ _0565_ _0007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2934_ _0024_ net61 net43 p_shaping_I.counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_1747_ _0793_ _0734_ _0723_ _0825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1678_ _0709_ _0662_ _0599_ _0756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1816_ _0793_ _0893_ _0894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2572__A1 _1363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2796_ _0280_ _0494_ _0495_ _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_13_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_55_Right_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_64_Right_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_66_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1601_ _0351_ _0676_ _0679_ _0680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_54_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1532_ _0609_ _0614_ _0615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2650_ _0334_ _0335_ _0338_ _0339_ _0341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_2581_ _0116_ _0267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_38_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input1_I BitIn vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1463_ _0036_ _0047_ _0058_ _0069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_1_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2015_ _1084_ _1085_ _1088_ _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2609__A2 _0049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2917_ _0013_ net59 clknet_1_1__leaf_CLK net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_2848_ _0527_ _0528_ _0551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2779_ _0415_ _0446_ _0449_ _0478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__1520__A2 _0602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1587__A2 _0663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_20_Left_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2702_ _0324_ _0323_ _0181_ _0381_ _0396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1515_ _0436_ _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2495_ _0167_ _0172_ _0173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2633_ _0284_ _0320_ _0321_ _0322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2564_ _0204_ _0033_ _0248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_10_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1446_ _1288_ _1299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_2_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_1_1__f_CLK clknet_0_CLK clknet_1_1__leaf_CLK vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_60_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2518__A1 _0051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output40_I net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2280_ _1353_ _1355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_51_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1799__A2 _0876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1995_ _1067_ _1069_ _1070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_42_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2616_ _0166_ _0266_ _0270_ _0304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2478_ _0059_ _0153_ _0154_ _0155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2547_ _1390_ _0229_ _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1899__I _0693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2935__D _0025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1780_ _0850_ _0857_ _0858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_12_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2332_ _1398_ _1405_ _1410_ _1411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_20_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2401_ _1433_ _0027_ _0071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2194_ _1261_ _1262_ _1263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2263_ _1321_ _1336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_35_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_23_Left_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1978_ _0719_ _1050_ _1051_ _1053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_30_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_51_Left_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_60_Left_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1832_ _0733_ _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1871__A1 _0542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1901_ _0739_ _0976_ _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2881_ _0578_ _0012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1763_ _0752_ _0840_ _0841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1694_ _0329_ _0709_ _0626_ _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_57_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2246_ _0124_ _1317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2315_ _1388_ _1391_ _1392_ _1393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1862__B2 _0770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2177_ _1214_ _1218_ _1246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_23_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput25 net25 Q[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput36 net52 addQ[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput14 net14 I[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_66_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1605__A1 _0318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2100_ _1090_ _0975_ _1171_ _0927_ _1172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_22_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2097__A1 _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2031_ _1104_ _1057_ _1105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_45_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_37_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1815_ _0708_ _0641_ _0648_ _0893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_43_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2933_ p_shaping_Q.bit_in_1 net62 net48 p_shaping_Q.bit_in_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2864_ Reg_Delay_Q.In net1 _0265_ _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2795_ _0063_ _0494_ _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1746_ _0797_ _0798_ _0824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2021__A1 _0666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1677_ _0711_ _0755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2229_ _1268_ _1298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_67_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2012__A1 _0739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1600_ _0677_ _0678_ _0679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1531_ _0611_ _0612_ _0613_ _0614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1462_ net32 _0058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2580_ _0210_ _0212_ _0264_ _0193_ _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_38_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2014_ _1085_ _1087_ _1084_ _1088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_9_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2916_ _0012_ net58 clknet_1_0__leaf_CLK net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2778_ _0453_ _0476_ _0477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2847_ _0529_ _0550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1729_ _0806_ _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_0_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_56_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2536__A2 _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2436__I _0108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2171__I _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2701_ _0100_ _0292_ _0293_ _0384_ _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_2632_ _0288_ _0294_ _0321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_6_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1514_ _0592_ _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_50_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1445_ net53 _1288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2494_ _0114_ _0112_ _0161_ _0167_ _0172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_2_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2563_ _0207_ _0247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_10_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2463__A1 _0096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2518__A2 _1403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2454__A1 _1367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout60 net65 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_67_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2693__B2 _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1994_ _1014_ _1018_ _1068_ _1069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2445__A1 _0051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2615_ _0271_ _0302_ _0303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2477_ _0140_ _0143_ _0137_ _0139_ _0154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2546_ _0217_ _0228_ _0229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_33_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1478__A2 _0080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2427__A1 _0096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2400_ _0066_ _0067_ _0068_ _0070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_12_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2902__A2 _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2331_ _1406_ _1301_ _1409_ _1279_ _1410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2262_ _1258_ _1335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_20_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2193_ _1236_ _1243_ _1260_ _1262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1977_ _1050_ _1051_ _0706_ _1052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_47_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2529_ _0199_ _0209_ _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_11_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2409__A1 _0077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1831_ _0840_ _0860_ _0752_ _0908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1900_ _0637_ _0975_ _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2880_ _0370_ _0576_ _0578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_32_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1693_ _0770_ _0771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1762_ _0839_ _0768_ _0840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2176_ _1243_ _1244_ _1245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2245_ _0200_ _1316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2314_ _1324_ _1386_ _1345_ _1392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__1523__I p_shaping_I.bit_in_1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput26 net26 Q[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput37 net51 addQ[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput15 net15 I[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_66_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2030_ _1044_ _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_57_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2932_ Reg_Delay_Q.Out net63 net47 p_shaping_Q.bit_in_1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_37_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2021__A2 _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1814_ _0479_ _0489_ _0691_ _0892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1745_ _0808_ _0815_ _0821_ _0822_ _0823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_2863_ _0611_ net42 _0564_ _0006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2794_ _0096_ _0273_ _0473_ _0375_ _0493_ _0494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_1676_ _0553_ _0754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_40_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1835__A2 _0911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2159_ _1126_ _0914_ _0712_ _1129_ _1228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__2793__B _1329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2228_ _1294_ _1296_ _1297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1461_ net55 _0047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1530_ p_shaping_I.ctl_1 _0612_ _0613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2013_ _0967_ _0732_ _1086_ _1087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_2915_ _0011_ net56 clknet_1_0__leaf_CLK net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_60_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1728_ _0673_ _0806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_33_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2846_ _0547_ _0548_ _0549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2777_ _0471_ _0475_ _0476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_5_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1659_ _0655_ _0683_ _0737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1808__A2 _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1983__A1 _1049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2700_ _0391_ _0136_ _0392_ _0394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2631_ _0292_ _0048_ _0049_ _0247_ _0320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_2_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2562_ _1277_ _1329_ _0246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_15_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1513_ net40 _0592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1444_ _1268_ _1277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2493_ _0171_ net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_61_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2829_ _0485_ _0508_ _0509_ _0531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_1_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2454__A2 _1403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1965__A1 _0887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout50 net39 net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout61 net64 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2445__A2 _0105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2693__A2 _1416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1993_ _0966_ _1013_ _1068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_15_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2545_ _0226_ _0227_ _0228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2614_ _0280_ _0301_ _0159_ _0302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2476_ _1397_ _0129_ _1281_ _0153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_65_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2216__B _0091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2192_ _1236_ _1243_ _1260_ _1261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2261_ _1280_ _1333_ _0211_ _1334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2330_ _1296_ _1313_ _1407_ _1349_ _1409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_55_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1976_ _0720_ _0755_ _1051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_43_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2528_ _0184_ _0201_ _0202_ _0206_ _0208_ _0209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_2459_ _1406_ _0129_ _0133_ _0134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_66_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_26_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1761_ _0585_ _0657_ _0667_ _0839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_1830_ _0862_ _0861_ _0902_ _0906_ _0907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_52_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1692_ _0569_ _0770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2313_ _1390_ _1391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_57_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2175_ _1238_ _1242_ _1244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2244_ _1311_ _1313_ _1314_ _1310_ _1315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_48_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2635__I _1406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1695__B _0636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1959_ _0883_ _0898_ _0939_ _0993_ _1034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_31_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput38 net38 addQ[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput27 net27 Q[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput16 net16 I[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_19_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2566__A1 _0100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2931_ _0002_ _2931_/E _2931_/RN p_shaping_Q.ctl_1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XFILLER_0_9_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1744_ _0656_ _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1813_ _0889_ _0890_ _0891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2862_ bit2symb.regi _0265_ _0564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2793_ _0492_ _1440_ _1329_ _1437_ _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_13_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1675_ _0752_ _0668_ _0753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1534__I p_shaping_Q.bit_in_1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2089_ _1161_ net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2158_ _1074_ _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2227_ _1295_ _1296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_39_Left_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_48_Left_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2476__S _1281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_57_Left_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1460_ net54 _0036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_66_Left_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_60_Right_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2012_ _0739_ _0854_ _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__2134__B _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2914_ _0010_ net57 clknet_1_0__leaf_CLK net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2845_ _0536_ _0537_ _0546_ _0548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_5_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1727_ _0705_ _0805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1658_ _0735_ _0714_ _0693_ _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_5_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2776_ _0233_ _0474_ _0611_ _0475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_13_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1589_ _0624_ _0657_ _0667_ _0668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_0_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1512_ _0569_ _0577_ _0393_ _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_54_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2492_ _0090_ _0170_ _0171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_2_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2561_ _0052_ _1439_ _0071_ _0221_ _0245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_2630_ _0316_ _0307_ _0317_ _0319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_49_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1443_ _1258_ _1268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_53_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2828_ _0485_ _0508_ _0530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_18_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2759_ _0283_ _0454_ _0455_ _1432_ _0426_ _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_TAPCELL_ROW_1_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout51 net37 net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout62 net64 net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_36_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2502__B _0039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1992_ _1022_ _1066_ _1067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_51_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2475_ _0030_ _0070_ _0081_ _0606_ _0152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__2381__A2 _1417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2544_ _0062_ _0145_ _0152_ _0227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2613_ _0281_ _0300_ _0301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_66_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1892__A1 _0818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1627__I _0542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1874__A1 _0942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2191_ _1235_ _1241_ _1259_ _1260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2260_ _1331_ _1291_ _1333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_47_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1975_ _0740_ _0742_ _0693_ _1050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__2051__A1 _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2527_ _1387_ _0207_ _0108_ _0208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_2458_ _0130_ _0132_ _0133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__1617__A1 _0694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2389_ _0053_ _0056_ _0046_ _0057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_34_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1760_ _0769_ _0835_ _0834_ _0838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1691_ _0753_ _0768_ _0769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_25_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2312_ _1389_ p_shaping_I.counter\[0\] _1390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_EDGE_ROW_27_Left_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2174_ _1238_ _1242_ _1243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2243_ _0069_ _1314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_11_Left_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2024__A1 _0844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput17 net17 Q[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_1889_ _0955_ _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput39 net39 addQ[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_1958_ _1030_ _1032_ _1033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xoutput28 net28 Q[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_31_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2600__B _0037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1688__S0 _0719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1796__B _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2930_ _0023_ net60 clknet_1_1__leaf_CLK bit2symb.regi vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2861_ _0563_ net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1743_ _0817_ _0819_ _0718_ _0820_ _0821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_1812_ _0869_ _0764_ _0890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1674_ Reg_Delay_Q.Out _0752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2792_ _0491_ _0176_ _0492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2226_ _1354_ _1295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2088_ _1158_ _1160_ _1161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2157_ _1226_ net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_63_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2291__I _1366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2011_ _0820_ _0916_ _0969_ _1085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_45_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2913_ _0009_ net56 clknet_1_0__leaf_CLK net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2844_ _0536_ _0537_ _0546_ _0547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1588_ _0658_ _0666_ _0553_ _0667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__1545__I _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1726_ p_shaping_Q.bit_in_2 _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1657_ _0457_ _0735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2775_ _0472_ _0473_ _0233_ _0474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2209_ _1276_ net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_56_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_14_Left_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1511_ _0532_ _0577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_50_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1442_ net54 _1258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2491_ _0093_ _0112_ _0169_ _0170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_2_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2560_ _0217_ _0228_ _0230_ _0242_ _0244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_65_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2696__A1 _0121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2758_ _1372_ _1293_ _1440_ _0455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2827_ _0527_ _0528_ _0529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_5_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1709_ _0785_ _0786_ _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2689_ _0059_ _0381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_1_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_1_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout52 net36 net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout63 net65 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_36_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2611__A1 _1329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2611__B2 _0184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1991_ _1033_ _1065_ _1066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2612_ _0283_ _0291_ net45 _0300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__2602__A1 _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2474_ _0145_ _0149_ _0608_ _0150_ _0151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2543_ _0148_ _0225_ _0226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_66_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1892__A2 _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout50_I net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1698__C _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_29_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1571__A1 _0647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2190_ _0942_ _1257_ _1149_ _0960_ _1259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_62_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1974_ _0688_ _0849_ _0989_ _1049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_47_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2823__A1 _0222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2339__B1 _1416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2526_ _1299_ _1369_ _0207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_2388_ _0054_ _1359_ _0055_ _0056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2457_ _0072_ _1296_ _0131_ _0132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_11_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2384__I _0051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1728__I _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_34_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1690_ _0754_ _0650_ _0757_ _0767_ _0768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XPHY_EDGE_ROW_2_Left_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2311_ p_shaping_I.counter\[1\] _1389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2242_ _1312_ _1313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_20_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2173_ _1241_ _1242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_63_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1957_ _0980_ _0982_ _1031_ _1032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_31_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1888_ _0964_ net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput29 net29 Q[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput18 net18 Q[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_2509_ _1320_ _1411_ _0188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1838__A2 _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2006__A2 _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1811_ _0425_ _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2791_ _0369_ _0491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2860_ _1396_ _0089_ _0563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_4_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1673_ _0731_ _0750_ _0725_ _0728_ _0668_ _0751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_1742_ _0806_ _0820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2190__A1 _0942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2225_ _1343_ _1294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2087_ _1115_ _1120_ _1159_ _1160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2156_ _1224_ _1225_ _1226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_36_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2010_ _0967_ _0631_ _0847_ _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2912_ _0008_ net63 clknet_1_1__leaf_CLK Reg_Delay_Q.Out vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_9_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1725_ _0789_ _0705_ _0724_ _0802_ _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_2843_ _0522_ _0525_ _0545_ _0546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2774_ _0097_ _0218_ _0248_ _0391_ _0462_ _0473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1656_ _0684_ _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_1587_ _0660_ _0663_ _0500_ _0665_ _0666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_0_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2702__A3 _0181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2208_ _0751_ _0836_ _1276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_56_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2139_ _1126_ _1051_ _1208_ _1209_ _1129_ _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_64_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1901__A1 _0739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2457__A2 _1296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1510_ net49 _0569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_2490_ _0114_ _0161_ _0167_ _0169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_61_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1708_ _0616_ _0750_ _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_41_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2826_ _0490_ _0507_ _0505_ _0528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2688_ _0193_ _0379_ _0380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_2757_ _0284_ _0078_ _0197_ _0454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1639_ _0382_ _0716_ _0717_ _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_1_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2387__I _1367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2439__A2 _0111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout64 net65 net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout42 net44 net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout53 net33 net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_20_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1990_ _0671_ _1063_ _1064_ _1065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_7_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2366__A1 _0031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2611_ _1329_ _1434_ _0295_ _0296_ _0184_ _0298_ _0299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai33_1
XFILLER_0_2_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2542_ _1383_ _0220_ _0223_ _1432_ _0224_ _0225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_2473_ _1385_ _0041_ _0060_ _0150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_2_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout43_I net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2809_ _0477_ _0481_ _0510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1874__A3 _0950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1973_ _1046_ _1047_ _0639_ _1048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_7_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2339__B2 _1417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2525_ _0203_ _0204_ _1285_ _0205_ _0206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_11_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2387_ _1367_ _0055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2456_ _0106_ _1366_ _0131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_11_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2511__A1 _0187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2776__S _0611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2502__A1 _1399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1654__I _0706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2172_ _1031_ _1131_ _1239_ _1240_ _1241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2310_ _1324_ _1345_ _1386_ _1388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2241_ _1258_ _1321_ _1312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_23_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1887_ _0907_ _0958_ _0963_ _0964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1956_ Reg_Delay_Q.Out _1031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_31_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1564__I net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput19 net19 Q[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2508_ _0059_ _0179_ _0183_ _0184_ _0186_ _0187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XTAP_TAPCELL_ROW_39_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2439_ _0095_ _0111_ _0112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2799__A1 _0440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1810_ _0631_ _0741_ _0816_ _0888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_57_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1741_ _0818_ _0714_ _0819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2790_ _0611_ _0438_ _0488_ _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1672_ _0732_ _0738_ _0744_ _0745_ _0749_ _0685_ _0750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_4
XANTENNA__1765__A2 _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2155_ _1168_ _1196_ _1198_ _1225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_36_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2224_ _1287_ _1290_ _1291_ _1292_ _1293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_63_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2086_ _1071_ _1112_ _1113_ _1159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_48_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1939_ _0956_ _0957_ _0907_ _1015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XOQPSK_PS_RCOSINE2_90 io_oeb[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_16_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1508__A2 _0542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1897__C _0754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1469__I net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_62_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1747__A2 _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_7_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1683__A1 _0647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2911_ _0007_ net60 clknet_1_1__leaf_CLK Reg_Delay_Q.In vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_EDGE_ROW_35_Left_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1724_ _0655_ _0794_ _0796_ _0799_ _0801_ _0802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_57_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_44_Left_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2842_ _0460_ _0544_ _0545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2773_ _0328_ _0330_ _0472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1655_ _0603_ _0733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1586_ _0664_ _0665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_0_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_53_Left_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2069_ _1109_ _1141_ _1142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2138_ _1126_ _0689_ _1209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2207_ _1269_ _1271_ _1275_ _1230_ _0960_ net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_28_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_64_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_62_Left_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1977__A2 _1051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_4_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2516__C _0101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1611__B _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2825_ _0523_ _0526_ _0527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_18_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_18_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1707_ _0771_ _0776_ _0784_ _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_53_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1638_ _0692_ _0678_ _0643_ _0717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_41_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2908__A1 _0234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2756_ _0437_ _0445_ _0435_ _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2687_ _0215_ _0214_ _0269_ _0341_ _0379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_1569_ _0371_ _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_39_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout65 net66 net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_36_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout54 net31 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout43 net44 net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2375__A2 _1337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2527__B _0108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1657__I _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2541_ _1309_ _0035_ _0224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2610_ _0054_ _0100_ _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2472_ _0148_ _0149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2437__B _0077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1567__I _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2808_ _0453_ _0476_ _0509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_41_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2739_ _0416_ _0433_ _0422_ _0435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_29_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2520__A2 _0044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1972_ _0819_ _0911_ _0743_ _1047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_55_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2339__A2 _1415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2524_ _0106_ _1358_ _0205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2455_ _1317_ _0130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_58_Right_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2386_ _1355_ _0054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_66_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_67_Right_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2018__A1 _0771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2018__B2 _0500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2569__A2 _0111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2171_ _0624_ _1240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2240_ _1289_ _1311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_7_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1886_ _0837_ _0904_ _0962_ _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1955_ _0685_ _1024_ _1028_ _1029_ _1030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_43_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_31_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2507_ _0185_ _0073_ _0103_ _0140_ _0186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2438_ _0099_ _0104_ _0110_ _0111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XTAP_TAPCELL_ROW_39_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2369_ _0032_ _0033_ _0034_ _0035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_34_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2723__A2 _1375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1671_ _0703_ _0747_ _0748_ _0749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1740_ _0629_ _0818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1665__I _0742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2085_ _1156_ _1157_ _1158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2154_ _1221_ _1223_ _1224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2223_ _0091_ _1292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2478__A1 _0059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XOQPSK_PS_RCOSINE2_80 io_oeb[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_33_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XOQPSK_PS_RCOSINE2_91 io_oeb[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_8_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1938_ _0966_ _1013_ _1014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_1869_ _0697_ _0910_ _0746_ _0946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_31_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2074__C _0771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2920__CLK clknet_1_0__leaf_CLK vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2880__A1 _0370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2249__C _0146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2910_ _0006_ net63 clknet_1_1__leaf_CLK p_shaping_I.bit_in vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_9_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2841_ _0159_ _0543_ _0544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1723_ _0603_ _0800_ _0801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1654_ _0706_ _0732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2772_ _0461_ _0470_ _0471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_5_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1910__A3 _0939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1585_ _0643_ _0664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2206_ _1274_ _1275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2068_ _1129_ _1135_ _1139_ _0875_ _1140_ _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_2137_ _0660_ _0663_ _0975_ _1134_ _1208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__2871__A1 _1399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1959__A3 _0939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2824_ _0525_ _0526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1706_ _0674_ _0777_ _0783_ _0723_ _0784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_1637_ net37 net36 _0716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_41_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2755_ _0452_ net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2686_ _0367_ _0377_ _0378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_18_Left_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1499_ _0447_ _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1568_ _0633_ _0647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_52_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout44 _0004_ net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout55 net30 net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_1_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout66 net3 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_9_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2471_ _0254_ _0147_ _0148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2540_ _1378_ _0103_ _0221_ _0223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_2_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2807_ _0490_ _0507_ _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2738_ _0416_ _0422_ _0433_ _0434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2669_ _0244_ _0357_ _0359_ _0360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_29_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2817__A1 _0025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1971_ _0646_ _1046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_55_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1795__A1 _0770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2385_ _0052_ _1314_ _0053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2523_ _1358_ _1303_ _0204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_11_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2454_ _1367_ _1403_ _1420_ _0129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
Xinput1 BitIn net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2448__B _0121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1488__I net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2569__A3 _0187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2170_ _1131_ _1073_ _1239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1954_ _0909_ _1029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1885_ _0838_ _0959_ _0961_ _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_43_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2368_ _1438_ _0034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_3_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2437_ _0105_ _0107_ _0077_ _0109_ _0110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2506_ _1349_ _0185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_39_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2299_ _1337_ _1375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_22_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1931__A1 _0771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2867__I _0566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2487__A2 _0127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_6_Left_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1670_ _0697_ _0748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2222_ _0157_ _0047_ _1291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_21_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2084_ _1154_ _1155_ _1124_ _1157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2153_ _1222_ _1223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XOQPSK_PS_RCOSINE2_92 io_oeb[32] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1937_ _0984_ _1012_ _1013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XOQPSK_PS_RCOSINE2_81 io_oeb[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_33_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XOQPSK_PS_RCOSINE2_70 io_oeb[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_8_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1868_ _0747_ _0944_ _0825_ _0945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1799_ _0875_ _0876_ _0877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_31_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1591__I _0669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1766__I _0308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2597__I _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1676__I _0553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2771_ _0267_ _0466_ _0469_ _0416_ _0470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2840_ _0063_ _0540_ _0541_ _0543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1722_ _0598_ _0684_ _0800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1653_ _0730_ _0731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1584_ _0662_ _0663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2699__A2 _1415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2205_ _1272_ _1273_ _1261_ _1274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_0_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2067_ _0718_ _1003_ _1140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_48_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2136_ _1073_ _1205_ _1206_ _1207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_fanout59_I net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1705_ _0742_ _0779_ _0780_ _0782_ _0783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__1959__A4 _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2754_ _0448_ _0451_ _0452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2823_ _0222_ _0367_ _0524_ _0146_ _0525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_1567_ _0645_ _0646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1636_ _0707_ _0710_ _0712_ _0714_ _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_2685_ _1318_ _0272_ _0373_ _0376_ _0377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_1498_ _0436_ _0447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2119_ _1075_ _0855_ _0602_ _1191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_1_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout56 net57 net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_44_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2470_ _0610_ _0613_ _0147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_23_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2806_ _0505_ _0506_ _0507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2737_ _0162_ _0432_ _0433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2668_ _0317_ _0358_ _0256_ _0359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_67_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1619_ _0457_ _0658_ _0697_ _0698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2599_ _0055_ _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_64_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2269__B1 _1340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1619__I0 _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1970_ _0873_ _0877_ _0945_ _0950_ _1045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_28_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2522_ _0076_ _0203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_11_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2453_ _0117_ _0127_ _0128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2384_ _0051_ _0052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput2 EN net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_34_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1594__I net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1701__A2 _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1884_ _0960_ _0902_ _0861_ _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1953_ _1025_ _1026_ _1027_ _1028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_28_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2505_ _1341_ _0184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_11_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_22_Left_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2459__B _0133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2436_ _0108_ _0109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2367_ _1433_ _1337_ _0033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_2298_ _1362_ _1374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_66_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1695__A1 _0720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2152_ _1200_ _1201_ _1220_ _1222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_2221_ _1289_ _1290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_17_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2083_ _1124_ _1154_ _1155_ _1156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1936_ _0671_ _1010_ _1011_ _1012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1867_ _0853_ _0943_ _0816_ _0944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XOQPSK_PS_RCOSINE2_93 io_oeb[33] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XOQPSK_PS_RCOSINE2_82 io_oeb[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XOQPSK_PS_RCOSINE2_71 io_oeb[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_58_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1798_ _0746_ _0765_ _0826_ _0876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_12_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2419_ _1396_ _0089_ _0090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_47_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1721_ _0797_ _0798_ _0799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1840__A1 _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2770_ _0466_ _0467_ _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1652_ _0702_ _0730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1583_ _0661_ _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_0_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2699__A3 _0033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2135_ _1031_ _1205_ _1206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2204_ _1236_ _1243_ _1260_ _1273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_48_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2066_ _0936_ _1138_ _1074_ _1139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_8_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1919_ _0985_ _0986_ _0994_ _0995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_44_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2139__A2 _1051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2899_ _1227_ _0590_ _0591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2378__A2 _0044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1813__A1 _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1704_ _0648_ _0781_ _0782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_38_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2753_ _0449_ _0450_ _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2684_ _0375_ _0325_ _0376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2369__A2 _0033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2822_ _0610_ _0222_ _0524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1497_ net50 _0436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1566_ _0641_ _0642_ _0644_ _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1635_ _0713_ _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2049_ _0925_ _1122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2118_ _0809_ _0970_ _1190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_52_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout57 net58 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_36_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2805_ _0497_ _0504_ _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1618_ _0318_ _0628_ _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_26_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2736_ _0423_ _0430_ _0431_ _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_14_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2667_ _0271_ _0302_ _0025_ _0358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1549_ _0627_ _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2598_ _0174_ _0284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_28_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2269__A1 _1337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2744__A2 _0203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2521_ _0039_ _1350_ _0043_ _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2383_ _1299_ _0051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2452_ _0118_ _0119_ _0122_ _0126_ _0127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput3 RST net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2680__A1 _0369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2719_ _0413_ net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2735__A2 _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1474__A2 net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1785__I p_shaping_Q.bit_in_1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2923__CLK clknet_1_0__leaf_CLK vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_63_Right_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_48_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1883_ _0669_ _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1952_ _0971_ _0854_ _0852_ _1027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_28_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2435_ _0135_ _1346_ _0108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_24_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2504_ _1294_ _0180_ _0181_ _1375_ _0182_ _0183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_47_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2366_ _0031_ _1368_ _0032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_2297_ _1357_ _1364_ _1370_ _1372_ _1373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_63_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1695__A2 _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2892__A1 _0844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2644__A1 _1357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2082_ _1150_ _1153_ _1133_ _1155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2151_ _1200_ _1201_ _1220_ _1221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2883__A1 _0203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2220_ _1430_ _1289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_48_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XOQPSK_PS_RCOSINE2_72 io_oeb[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1935_ _0701_ _1009_ _0995_ _0996_ _1011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_56_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1797_ _0603_ _0874_ _0875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1866_ _0687_ _0713_ _0943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XOQPSK_PS_RCOSINE2_94 io_oeb[34] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XOQPSK_PS_RCOSINE2_83 io_oeb[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2418_ _1413_ _0088_ _0089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2349_ _1347_ _1429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_66_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1601__A2 _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_7_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1651_ _0729_ net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_65_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1720_ _0425_ _0713_ _0798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_41_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1582_ net51 net52 _0661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_0_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1659__A2 _0683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2065_ _0928_ _1137_ _1138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2203_ _1245_ _1247_ _1272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2134_ _1202_ _1204_ _0624_ _1131_ _1205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_44_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1883__I _0669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1918_ _0993_ _0994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1849_ _0351_ _0866_ _0926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2898_ _0582_ _0589_ _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_4_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2821_ _0518_ _0522_ _0523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_14_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1703_ _0716_ _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1634_ _0651_ _0640_ _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_30_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2683_ _0374_ _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2752_ _0407_ _0412_ _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1565_ _0643_ _0644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_1496_ _0340_ _0414_ _0425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_1_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2048_ _1121_ net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2117_ _0562_ _0624_ _0604_ _1189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA_fanout64_I net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout58 net59 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout47 _0005_ net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_36_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2532__A3 _0127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_41_Left_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_50_Left_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_66_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2804_ _0497_ _0504_ _0505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1617_ _0694_ _0695_ _0696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1970__A1 _0873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2597_ _0282_ _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_1_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2666_ _0114_ _0025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2735_ _1428_ _0430_ _0431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1722__A1 _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1548_ net38 _0627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1479_ _1397_ _0233_ _0243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_49_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2450__A2 _0048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2451_ _0108_ _1415_ _0123_ _0125_ _0126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_2520_ _1351_ _0044_ _0101_ _0027_ _0201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_36_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2382_ _0046_ _0048_ _0049_ _0050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_52_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2680__A2 _0176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2718_ _0407_ _0412_ _0413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2499__A2 _0176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2649_ _0168_ _1377_ _1370_ _1406_ _0339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_37_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1882_ _0862_ _0861_ _0902_ _0959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1951_ _0817_ _0631_ _0636_ _0976_ _1026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_24_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2365_ _1430_ _0031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_3_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2503_ _1356_ _1375_ _0182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2434_ _0106_ _1343_ _1441_ _1438_ _0107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_2296_ _1371_ _1372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_63_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2405__A2 _0048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2341__A1 _1301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2644__A2 _1364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1907__A1 _0752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2081_ _1133_ _1150_ _1153_ _1154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_2150_ _1207_ _1219_ _1220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2883__A2 _1422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1934_ _0701_ _0995_ _0996_ _1009_ _1010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_56_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XOQPSK_PS_RCOSINE2_73 io_oeb[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_29_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XOQPSK_PS_RCOSINE2_84 io_oeb[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1796_ _0810_ _0777_ _0673_ _0874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1865_ _0605_ _0879_ _0942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_3_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XOQPSK_PS_RCOSINE2_95 io_oeb[35] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2874__A2 _0176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2417_ _1391_ _0083_ _0087_ _0088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2348_ _0607_ _1428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2571__A1 _0252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2913__CLK clknet_1_0__leaf_CLK vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2279_ _0036_ _1353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_50_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2562__A1 _1277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1650_ _0668_ _0728_ _0729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1581_ _0659_ _0660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_13_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2202_ _1222_ _1248_ _1251_ _1270_ _1271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_28_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2064_ _0809_ _1136_ _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2133_ _1203_ _1204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_63_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1917_ _0887_ _0987_ _0992_ _0758_ _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_2897_ _0582_ _0775_ _0566_ _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_29_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1848_ _0788_ _0925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1779_ _0852_ _0853_ _0856_ _0857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_12_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2820_ _0267_ _0519_ _0520_ _0416_ _0522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_2751_ _0366_ _0406_ _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1702_ _0329_ _0626_ _0629_ _0542_ _0780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_53_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1564_ net50 _0643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1633_ _0664_ _0711_ _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_41_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2682_ _0282_ _0374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1495_ net38 _0414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2047_ _1115_ _1120_ _1121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2116_ _1178_ _1187_ _1188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_9_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout59 net66 net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout48 _0005_ net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2765__A1 _0273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1843__B _0706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2517__A1 _0031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1559__A2 _0636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2508__B2 _0184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2508__A1 _0059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2444__B1 _1415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2803_ _0267_ _0502_ _0503_ _0234_ _0504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2734_ _0208_ _0424_ _0427_ _0184_ _0429_ _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_14_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1722__A2 _0684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1616_ _0521_ _0592_ _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1663__B _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1547_ _0625_ _0626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2596_ _1383_ _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2665_ _0316_ _0303_ _0307_ _0357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1478_ _1419_ _0080_ _0146_ _0222_ _0233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_37_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1477__A1 _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2450_ _1326_ _0048_ _0125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_23_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2381_ _1402_ _1417_ _1401_ _0049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_11_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2717_ _0310_ _0408_ _0411_ _0412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_65_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2648_ _0046_ _0337_ _1383_ _0338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_10_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2579_ _0258_ _0261_ _0263_ _0264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_25_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2187__A2 _0754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2111__A2 _1051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1870__A1 _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1950_ _0852_ _1025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1478__B _0146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1881_ _0956_ _0957_ _0958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1925__A2 _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2502_ _1399_ _1311_ _0039_ _0181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_2433_ _0157_ _0106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2364_ _1432_ _1435_ _0026_ _0029_ _0030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__2350__A2 _1429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2295_ _1408_ _1371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_59_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2405__A3 _0049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1852__A1 _0927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2238__I _0091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2080_ _0731_ _1151_ _1152_ _0672_ _1153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__2096__A1 _0731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XOQPSK_PS_RCOSINE2_85 io_oeb[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XOQPSK_PS_RCOSINE2_96 io_oeb[36] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1933_ _0998_ _1008_ _1009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_44_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_26_Left_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XOQPSK_PS_RCOSINE2_74 io_oeb[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_8_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1864_ _0939_ _0940_ _0941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1795_ _0770_ _0868_ _0872_ _0873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_3_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2347_ _1414_ _1426_ _1427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2416_ _0084_ _0085_ _0086_ _1389_ _0087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2278_ _1349_ _1309_ _1351_ _1352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_10_Left_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2933__D p_shaping_Q.bit_in_1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2562__A2 _1329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1580_ _0489_ _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2132_ _0889_ _0511_ _1203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2201_ _1263_ _1270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2063_ _0660_ _0714_ _1136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1847_ _0908_ _0923_ _0924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_60_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1916_ _0806_ _0935_ _0988_ _0991_ _0992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_2896_ _1038_ _0774_ _0586_ _0570_ _0809_ _0018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__2792__A2 _0176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1778_ _0854_ _0855_ _0665_ _0856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1701_ _0778_ _0676_ _0779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_53_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2750_ _0415_ _0446_ _0448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_2681_ _0368_ _0247_ _0372_ _0373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1494_ _0308_ _0393_ _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1563_ _0371_ _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1632_ _0651_ _0675_ _0414_ _0711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_1_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2526__A2 _1369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2115_ _0730_ _1186_ _1187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XOQPSK_PS_RCOSINE2_100 io_oeb[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xfanout49 net41 net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_64_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2046_ _1116_ _1119_ _1120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_57_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2879_ _0491_ _0574_ _0576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_13_Left_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2692__A1 _0105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2444__A1 _1314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2444__B2 _0101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2802_ _0380_ _0502_ _0503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2664_ _0319_ _0355_ _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2733_ _0132_ _0428_ _0282_ _0429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1615_ _0691_ _0661_ _0693_ _0694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_1546_ _0286_ _0625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_1477_ _0168_ _0189_ _0211_ _0222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_2595_ _0150_ _0156_ _0225_ _0608_ _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_1_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2029_ _1056_ _1102_ _1103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_45_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2380_ _1282_ _0058_ _0048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_23_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2647_ _1374_ _1407_ _0336_ _0337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2716_ _0360_ _0409_ _0410_ _0411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1529_ net63 _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2578_ _1279_ _1370_ _0262_ _0263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_25_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2895__A1 _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1880_ _0862_ _0954_ _0955_ _0924_ _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__1870__A2 _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_38_Left_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1478__C _0222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_47_Left_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2501_ _1416_ _0180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_39_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2432_ _1376_ _1302_ _0105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2363_ _1371_ _0028_ _1316_ _0029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2294_ _1367_ _1368_ _1369_ _1370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__1513__I net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_56_Left_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2102__A3 _0933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2638__A1 _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_65_Left_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_62_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1852__A2 _0928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1843__A2 _0663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XOQPSK_PS_RCOSINE2_97 io_oeb[37] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1863_ _0884_ _0899_ p_shaping_Q.bit_in_2 _0940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_56_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1932_ _0828_ _1001_ _1007_ _0880_ _1008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_44_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XOQPSK_PS_RCOSINE2_86 io_oeb[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XOQPSK_PS_RCOSINE2_75 io_oeb[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1794_ _0870_ _0871_ _0851_ _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__1952__B _0852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2415_ _1414_ _1426_ _0086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_24_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1531__A1 _0611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2346_ _1425_ _1426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2277_ _1350_ _1351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_66_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1589__A1 _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1761__A1 _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2062_ _0826_ _1023_ _0911_ _1134_ _0974_ _1135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_2200_ _1266_ _1267_ _1269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2131_ _1125_ _1202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_28_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2864__I1 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1846_ _0909_ _0918_ _0922_ _0923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_56_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1915_ _0867_ _0849_ _0989_ _0990_ _0851_ _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_1777_ _0790_ _0764_ _0855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2895_ _0763_ _0755_ _0587_ _0572_ _1075_ _0017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_8_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1504__A1 _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2329_ _1338_ _1407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_47_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1700_ _0628_ _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_53_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1631_ _0708_ _0709_ _0641_ _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_38_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2680_ _0369_ _0176_ _0113_ _0370_ _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_5_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1493_ _0329_ _0351_ _0382_ _0393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_1562_ _0640_ _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_1_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2045_ _1068_ _1117_ _1118_ _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_55_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2114_ _1179_ _1183_ _1185_ _1186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XOQPSK_PS_RCOSINE2_101 io_oeb[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_57_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1829_ _0882_ _0901_ _0906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2878_ _0575_ _0011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_9_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2453__A2 _0127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1587__B _0500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2692__A2 _0221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2801_ _0498_ _0501_ _0502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_14_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1707__A1 _0771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1970__A4 _0950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1955__A1 _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1614_ _0692_ _0371_ _0693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_41_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2594_ _0279_ _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2663_ _0332_ _0354_ _0355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2732_ _0131_ _1327_ _0174_ _0428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1545_ _0585_ _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_66_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1960__B _0694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2132__A1 _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1476_ _0200_ _0211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_22_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2028_ _1079_ _1096_ _1099_ _1101_ _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1946__A1 _0672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_20_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2646_ _0034_ _0203_ _0336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2715_ _0319_ _0355_ _0410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2577_ _1363_ _0195_ _0262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2916__CLK clknet_1_0__leaf_CLK vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1459_ _1430_ _1441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1528_ _0610_ _0611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_45_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2895__A2 _0755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2431_ _0100_ _0078_ _0103_ _1318_ _0104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2500_ _0174_ _0132_ _0177_ _0179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_39_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2293_ _1335_ _1365_ _1369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_2362_ _1292_ _0027_ _1439_ _1380_ _0028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__2638__A2 _1429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2629_ _0304_ _0306_ _0317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_0_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XOQPSK_PS_RCOSINE2_76 io_oeb[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1862_ _0886_ _0930_ _0938_ _0770_ _0939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_1793_ _0308_ _0720_ _0679_ _0871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_1931_ _0771_ _1006_ _1007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_33_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XOQPSK_PS_RCOSINE2_98 io_oeb[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XOQPSK_PS_RCOSINE2_87 io_oeb[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_3_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2414_ _0062_ _1386_ _0070_ _0081_ _0085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_2345_ _1348_ _1418_ _1421_ _1424_ _1425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_2276_ _0036_ _1430_ _1350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2547__A1 _1390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_41_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2130_ _1188_ _1195_ _1201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2061_ _1090_ _1134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_28_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1914_ _0308_ _0760_ _0869_ _0990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1845_ _0656_ _0921_ _0922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1776_ _0760_ _0854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2894_ _0647_ _0572_ _0663_ _0587_ _0016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_29_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2529__A1 _0199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1504__A2 _0500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2328_ _1404_ _1406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2701__A1 _0100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2259_ _0178_ _1331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1630_ _0628_ _0709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_53_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1492_ _0371_ _0382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_1561_ _0286_ _0640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XOQPSK_PS_RCOSINE2_102 io_oeb[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_2044_ _1020_ _1021_ _1066_ _1118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2113_ _1179_ _1184_ _1183_ _1185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_52_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2119__B _0602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2877_ _0491_ _0574_ _0575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2462__A3 _1369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1828_ _0905_ net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1759_ _0751_ _0836_ _0837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1725__A2 _0705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1622__I p_shaping_Q.counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2800_ _0374_ _0499_ _0501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2731_ _0285_ _0044_ _0426_ _0427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_14_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1613_ _0632_ _0692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1544_ _0623_ net47 _1544_/ZN vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2662_ _1391_ _0347_ _0353_ _0354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2593_ _0155_ _0225_ _0278_ _0607_ _0279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_66_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1475_ net35 _0200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1643__A1 _0719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2027_ _1029_ net46 _1101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_60_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2929_ p_shaping_I.bit_in_1 net65 net42 p_shaping_I.bit_in_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_20_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1928__A2 _0636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2714_ _0319_ _0355_ _0409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1527_ p_shaping_I.bit_in _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_2645_ _0109_ _0181_ _0335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2576_ _1279_ _0259_ _0260_ _0130_ _0261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__1864__A1 _0939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1458_ net32 _1430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_60_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2335__A2 _1330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2361_ _1291_ _0027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2430_ _0101_ _1340_ _0103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_39_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2292_ _1325_ _1368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_63_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2559_ _0191_ _0242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2628_ _0256_ _0316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1837__A1 _0742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1688__I1 _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2037__B _0672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2565__A2 _1361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1930_ _0842_ _1002_ _1003_ _1004_ _1005_ _1006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_TAPCELL_ROW_44_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XOQPSK_PS_RCOSINE2_88 io_oeb[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XOQPSK_PS_RCOSINE2_77 io_oeb[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1861_ _0931_ _0934_ _0937_ _0938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_56_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1792_ _0869_ _0764_ _0664_ _0778_ _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XOQPSK_PS_RCOSINE2_99 io_oeb[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_3_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2344_ _1278_ _1423_ _1424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2413_ _1428_ _0030_ _0041_ _0060_ _0084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2275_ _1308_ _1349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_47_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1625__I _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2060_ _1073_ _1132_ _1133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_44_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1913_ _0681_ _0709_ _0644_ _0989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_2893_ _0844_ _0587_ _0588_ _0015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1844_ _0919_ _0920_ _0404_ _0921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1775_ _0760_ _0662_ _0853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2327_ _1314_ _0113_ _1400_ _1403_ _1404_ _1363_ _1405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_2258_ _1327_ _1328_ _1329_ _1330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__2794__C _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2189_ _1109_ _1255_ _1256_ _1257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_26_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1873__C _0770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1560_ _0577_ _0639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_53_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XOQPSK_PS_RCOSINE2_103 io_oeb[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_2112_ _1001_ _1034_ _1041_ _1184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1491_ _0361_ _0371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_39_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2043_ _1020_ _1021_ _1066_ _1117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_52_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1827_ _0837_ _0904_ _0905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_60_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2876_ net2 _1361_ _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1758_ _0769_ _0835_ _0836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1725__A3 _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1689_ _0758_ _0766_ _0767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2730_ _0262_ _0323_ _0426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2661_ _1324_ _0348_ _0349_ _0350_ _0352_ _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_1612_ net50 _0691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1543_ _0623_ net42 _1543_/ZN vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1474_ _0178_ net34 _0189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_22_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2592_ _1398_ _0276_ _0277_ _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_66_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2026_ _0820_ _0782_ _0989_ _1097_ _1098_ _0893_ _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai33_1
XFILLER_0_15_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2928_ p_shaping_I.bit_in net61 net42 p_shaping_I.bit_in_1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2859_ _0557_ _0559_ _0561_ _0516_ _0232_ net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XPHY_EDGE_ROW_17_Left_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2371__A3 _0037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2362__A3 _1439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2464__I _0108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2644_ _1357_ _1364_ _0334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2713_ _0173_ _0231_ _0313_ _0356_ _0408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__2889__A1 _0486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1526_ _0243_ _0609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1457_ net35 _1408_ _1419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_10_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2575_ _1355_ _0194_ _0136_ _0051_ _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_2009_ _1034_ _1041_ _0789_ _1083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_9_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2549__I _1390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1855__A2 _0687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2360_ _1436_ _1437_ _1440_ _1368_ _1404_ _0026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_2291_ _1366_ _1367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_63_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2099__A2 _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_47_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2627_ _0315_ net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_56_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1509_ _0425_ _0511_ _0553_ _0562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XPHY_EDGE_ROW_34_Left_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2489_ _0163_ _0164_ _0165_ _0166_ _0167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_2558_ _0241_ net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1837__A2 _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_43_Left_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_53_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_52_Left_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1786__C _0700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XOQPSK_PS_RCOSINE2_67 io_oeb[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_56_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1860_ _0792_ _0895_ _0936_ _0719_ _0937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_44_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XOQPSK_PS_RCOSINE2_78 io_oeb[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XOQPSK_PS_RCOSINE2_89 io_oeb[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1791_ _0634_ _0869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2274_ _1346_ _1347_ _1316_ _1348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_2343_ _1422_ _1325_ _1423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2412_ _1323_ _1427_ _0061_ _0082_ _0083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__1977__B _0706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1989_ _0702_ _1042_ _1043_ _1062_ _1064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_TAPCELL_ROW_41_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1746__A1 _0797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_5_Left_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_6_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1843_ _0646_ _0663_ _0706_ _0920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1912_ _0816_ _0855_ _0988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2892_ _0844_ _0583_ _0588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1774_ _0851_ _0852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_52_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2257_ _0211_ _1408_ _1329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_2326_ _1346_ _1404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_55_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2188_ _0618_ _1255_ _1256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2465__A2 _0031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1976__A1 _0720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_31_Left_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2456__A2 _1366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2292__I _1325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1490_ net38 _0361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_53_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2042_ _1015_ _1014_ _1017_ _1067_ _1116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_55_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2111_ _0974_ _1051_ _1181_ _1182_ _1183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XOQPSK_PS_RCOSINE2_104 io_oeb[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_TAPCELL_ROW_52_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_17_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1826_ _0838_ _0861_ _0903_ _0904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XTAP_TAPCELL_ROW_60_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2875_ _1277_ _0572_ net44 _0573_ _0010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_13_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1757_ _0670_ _0833_ _0834_ _0835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1688_ _0761_ _0763_ _0765_ _0688_ _0719_ _0735_ _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_40_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2919__CLK clknet_1_0__leaf_CLK vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2309_ _1385_ _1386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2610__A2 _0100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_57_Right_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1456__I net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_66_Right_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1611_ _0687_ _0688_ _0689_ _0690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__2062__B1 _0911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2660_ _0149_ _0280_ _0352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1542_ _0612_ _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1473_ net53 _0178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2591_ _0175_ _0045_ _1318_ _0277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_65_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2025_ _0893_ _1097_ _1098_ _1099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input2_I EN vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2927_ _0000_ _2927_/E _2927_/RN p_shaping_I.ctl_1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XFILLER_0_9_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1809_ _0886_ _0887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_31_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2858_ _0551_ _0560_ _0547_ _0561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2789_ _0146_ _0222_ _0487_ _0488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_13_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2108__A1 _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2822__A2 _0222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2712_ _0366_ _0406_ _0407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_2574_ _0107_ _0142_ _0259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2643_ _0210_ _0212_ _0264_ _0192_ _0333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_1456_ net34 _1408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_1525_ _0607_ _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_10_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2008_ _1073_ _1081_ _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_fanout60_I net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2577__A1 _1363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output41_I net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1607__A3 _0683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2568__A1 _0096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2290_ _0178_ _1366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_63_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_47_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2557_ _0173_ _0231_ _0240_ _0241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2626_ _0310_ _0314_ _0315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1508_ _0521_ _0542_ _0553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_49_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2488_ _1389_ _0166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2798__A1 _0080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1470__A1 _0091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2722__A1 _0369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1790_ _0795_ _0866_ _0867_ _0848_ _0577_ _0868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_56_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XOQPSK_PS_RCOSINE2_79 io_oeb[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2789__A1 _0146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XOQPSK_PS_RCOSINE2_68 io_oeb[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2244__B _1314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2411_ _0063_ _1386_ _0070_ _0081_ _0082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2342_ _0189_ _1422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2273_ _0036_ _0047_ net33 _0058_ _1347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
X_1988_ _0702_ _1042_ _1043_ _1062_ _1063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_47_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2609_ _0292_ _0049_ _0296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_65_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1746__A2 _0798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1773_ _0592_ _0851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1911_ _0694_ _0756_ _0987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1842_ _0665_ _0649_ _0781_ _0919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_44_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1737__A2 _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2891_ _0586_ _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2187_ _1134_ _0754_ _1254_ _1202_ _1255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_2256_ _1300_ _1291_ _1299_ _1328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2325_ _1379_ _1401_ _1402_ _1403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__1673__A1 _0731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1976__A2 _0755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2041_ _1071_ _1114_ _1115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2110_ _0808_ _1137_ _1029_ _1182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_60_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1825_ _0862_ _0902_ _0903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1756_ _0787_ _0832_ _0834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2080__A1 _0731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2874_ _0570_ _0176_ _0573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1687_ _0764_ _0642_ _0708_ _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2308_ _1348_ _1352_ _1373_ _1384_ _1385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_0_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1646__A1 _0705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2393__I p_shaping_I.bit_in_1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2239_ _1306_ _1307_ _1308_ _1309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_0_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2062__A1 _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1610_ _0635_ _0652_ _0682_ _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_41_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2590_ _0272_ _0274_ _0275_ _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_66_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2117__A2 _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1541_ _0618_ net47 _0622_ _0002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1472_ _0157_ _1365_ _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_22_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2024_ _0844_ _0971_ _1075_ _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__1800__A1 _0873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2926_ _0022_ net62 net48 p_shaping_Q.counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2857_ _0536_ _0537_ _0546_ _0560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_9_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1808_ _0569_ _0598_ _0886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1739_ _0816_ _0817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2788_ _0486_ _0080_ _0487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_54_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2711_ _0378_ _0405_ _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_50_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1524_ _0606_ _0607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2573_ _0140_ _0257_ _0258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2642_ _0328_ _0331_ _0332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2001__I _0818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1455_ _1277_ _1310_ _1387_ _1397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_10_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2510__A2 _0111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2007_ _0887_ _1049_ _1077_ _1080_ _1081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_25_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2909_ _0025_ _0597_ _0024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output34_I net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_0_CLK CLK clknet_0_CLK vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_24_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1507_ _0532_ _0542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2487_ _0117_ _0127_ _0165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_23_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2556_ _0090_ _0170_ _0239_ _0240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__2731__A2 _0044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2625_ _0173_ _0231_ _0313_ _0314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_38_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2798__A2 _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2722__A2 _1361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2789__A2 _0222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XOQPSK_PS_RCOSINE2_69 io_oeb[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_44_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2525__B _1285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1655__I _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2341_ _1301_ _1420_ _1280_ _1421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_24_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2410_ _0074_ _0075_ _0079_ _1382_ _0081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_2272_ _0124_ _1346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_20_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1987_ _1044_ _1057_ _1060_ _1061_ _1062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_15_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2539_ _0125_ _0221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2608_ _0054_ _0294_ _0295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_58_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2640__A1 _0252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2080__B _0672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1475__I net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2459__A1 _1406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1910_ _0884_ _0899_ _0939_ _0986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_44_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2890_ _0582_ _0567_ _0586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1841_ _0843_ _0912_ _0917_ _0852_ _0918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1772_ _0637_ _0763_ _0847_ _0849_ _0639_ _0850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_40_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2324_ _1305_ _1402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2186_ _1134_ _0968_ _1227_ _1254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2255_ _1441_ _1325_ _0102_ _1326_ _1327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_63_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1509__B _0553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2040_ _1112_ _1113_ _1114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_60_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2873_ _0570_ _0572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_17_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1755_ _0787_ _0832_ _0833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1824_ _0882_ _0901_ _0902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1686_ _0640_ _0764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_0_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2238_ _0091_ _1308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2307_ _1377_ _1381_ _1383_ _1384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1646__A2 _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2169_ _1236_ _1237_ _1238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_0_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1702__B _0542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1540_ net47 _0621_ _0622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_22_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1471_ net54 _0157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_65_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2023_ _0807_ _0969_ _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1807_ _0804_ _0884_ _0885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_57_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2925_ _0021_ net61 net48 p_shaping_Q.counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2856_ _0530_ _0533_ _0558_ _0559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1738_ _0599_ _0816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1669_ _0647_ _0659_ _0746_ _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_40_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2787_ _0374_ _0486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_36_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_31_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2504__B1 _0181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2710_ _0114_ _0402_ _0403_ _0405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__1607__B _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1523_ p_shaping_I.bit_in_1 _0606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2572_ _1363_ _1360_ _0247_ _0257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2641_ _0094_ _0330_ _0331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1454_ _1343_ _1376_ _1387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_65_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2006_ _1078_ _0889_ _1079_ _1080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2026__A2 _0782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2908_ _0234_ p_shaping_I.counter\[0\] _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2839_ _0280_ _0540_ _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2017__A2 _0754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2258__B _1329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1767__A1 _0844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2624_ _0311_ _0312_ _0240_ _0313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_6_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1506_ net40 _0532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2555_ _0093_ _0172_ _0238_ _0239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2486_ _0156_ _0162_ _0152_ _0164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_2_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2682__I _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_24_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1921__A1 _0873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2271_ _1344_ _1345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2340_ _1376_ _1312_ _1331_ _1420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_20_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2477__A2 _0143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1986_ _1044_ _1055_ _1061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2607_ _0292_ _0293_ _0294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_11_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1581__I _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2538_ _0218_ _0195_ _0219_ _1374_ _1378_ _0220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_2469_ _1398_ _0134_ _0137_ _0139_ _0144_ _0145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__2468__A2 _0143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1979__A1 _1049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1840_ _0813_ _0913_ _0915_ _0916_ _0917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_56_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2631__A2 _0048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1771_ _0848_ _0849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2395__A1 _1296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2254_ _0178_ _1326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2323_ _1283_ _1401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_20_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2497__I _1285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2185_ _1253_ net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_63_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1969_ _0880_ _1044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_9_Left_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_53_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2392__A4 _0060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2803__C _0234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2129__A1 _0731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1823_ _0885_ _0899_ _0900_ _0901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_60_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2872_ _0571_ _0009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2604__A2 _1429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1754_ _0788_ _0803_ _0831_ _0832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_52_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1685_ _0762_ _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2306_ _1382_ _1383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2237_ _1283_ _1307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_0_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2099_ _0967_ _0813_ _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_51_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2168_ _1232_ _1235_ _1237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_0_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_8_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1470_ _0091_ _0113_ _0124_ _0135_ _0146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_1_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_65_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_59_Left_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2022_ _0666_ _0710_ _1095_ _1096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2589__A1 _1281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1806_ _0883_ _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2924_ _0020_ net60 clknet_1_1__leaf_CLK net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2786_ _0484_ _0485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2855_ _0529_ _0549_ _0558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_62_Right_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1599_ _0361_ _0678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1668_ _0682_ _0746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1737_ _0809_ _0811_ _0814_ _0815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_40_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2504__B2 _1375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2036__S _0942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2640_ _0252_ _0253_ _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1522_ _0605_ _0005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1453_ _1365_ _1376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_22_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2571_ _0252_ _0255_ _0256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2005_ _0822_ _1079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2907_ _0596_ _0023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1584__I _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2734__B2 _0184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2769_ _0291_ _0379_ _0193_ _0467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2838_ _0538_ _0539_ _0540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2554_ _0232_ _0235_ _0236_ _0237_ _0238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_2_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2623_ _0242_ _0230_ _0312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1505_ net49 _0521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2485_ _0152_ _0156_ _0162_ _0163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1455__A1 _1277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1749__A2 _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2270_ _1330_ _1334_ _1342_ _1344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_59_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1985_ _0863_ _0997_ _1059_ _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2732__B _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2606_ _1356_ _0293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_2_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2537_ _1351_ _0044_ _0219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2399_ _1382_ _0040_ _0068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2468_ _0140_ _0143_ _0144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_38_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2476__I0 _1397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1705__C _0782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1667__A1 _0694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1770_ _0677_ _0625_ _0759_ _0447_ _0848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_37_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2631__A3 _0049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2184_ _1248_ _1252_ _1253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2322_ _1277_ _1399_ _1400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2253_ net31 net30 _1325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_20_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_40_Left_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2446__C _0031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_25_Left_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1968_ _0985_ _1034_ _1041_ _1043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1899_ _0693_ _0975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1897__B2 _0791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2138__A2 _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1649__A1 _0672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2598__I _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2065__A1 _0928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1822_ _0804_ _0884_ _0899_ _0788_ _0900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_TAPCELL_ROW_60_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1753_ _0804_ _0805_ _0823_ _0830_ _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2871_ _1399_ _0570_ _0571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_25_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1879__A1 _0669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1684_ _0677_ _0297_ _0600_ _0762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_20_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2167_ _1232_ _1235_ _1236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2305_ _0135_ _1382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2236_ _1305_ _1306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2098_ _1090_ _1025_ _0932_ _1170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_51_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2359__A2 _1439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2906__I1 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1497__I net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2021_ _0666_ _0710_ _1025_ _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2923_ _0019_ net58 clknet_1_0__leaf_CLK net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XANTENNA__2791__I _0369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1805_ _0705_ _0724_ _0802_ _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_53_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1736_ _0812_ _0813_ _0755_ _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_2785_ _0471_ _0475_ _0483_ _0484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2854_ _0555_ _0556_ _0557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1667_ _0694_ _0695_ _0745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1598_ _0632_ _0677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2219_ _1286_ _1287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_63_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_12_Left_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2570_ _0094_ _0253_ _0255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1521_ _0404_ _0562_ _0585_ _0604_ _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_1452_ _1354_ _1365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2004_ _0974_ _1078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_45_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_33_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2906_ bit2symb.regi net1 _0595_ _0596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2431__A1 _0100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1719_ _0708_ _0641_ _0644_ _0648_ _0797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_26_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2699_ _0324_ _1415_ _0033_ _0392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2768_ _0381_ _0464_ _0465_ _0466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_2837_ _0370_ _0462_ _0486_ _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2413__B2 _0060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1504_ _0457_ _0500_ _0511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2922__CLK clknet_1_0__leaf_CLK vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2553_ _0112_ _0237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2622_ _0167_ _0172_ _0311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2484_ _0158_ _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_58_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_38_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2327__S1 _1363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1595__I _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_0_CLK_I CLK vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2882__A1 _0370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1984_ _1058_ _1048_ _0822_ _1059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_23_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2929__RN net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2605_ _0052_ _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2467_ _0034_ _0141_ _0107_ _0142_ _0143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_2536_ _1310_ _0168_ _0218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_2398_ _1371_ _0032_ _0037_ _0067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_3_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2321_ _1286_ _1399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2183_ _1222_ _1251_ _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2252_ _1323_ _1324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_63_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1967_ _0985_ _1034_ _1041_ _1042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1898_ _0732_ _0974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_43_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2519_ _0121_ _0196_ _0198_ _0199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_54_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2837__A1 _0370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2870_ net2 _0570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_17_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1693__I _0770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1821_ _0898_ _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1752_ _0824_ _0825_ _0827_ _0829_ _0830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_52_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1683_ _0647_ _0760_ _0761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2304_ _1378_ _1380_ _1381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2540__A3 _0221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1642__B _0720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2097_ _0826_ _1023_ _0801_ _1169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_45_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2166_ _1179_ _1233_ _1234_ _1122_ _1235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_2235_ _1268_ _1305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_0_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_51_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_66_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2020_ _1044_ _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_57_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1797__A1 _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2922_ _0018_ net58 clknet_1_0__leaf_CLK net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__2589__A3 _0273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2853_ _0526_ _0545_ _0522_ _0556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1666_ _0660_ _0653_ _0741_ _0743_ _0744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_1804_ _0865_ _0881_ _0882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1735_ _0676_ _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2784_ _0461_ _0470_ _0483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_13_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1721__A1 _0797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1597_ _0651_ _0675_ _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2149_ _1214_ _1218_ _1219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_36_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2218_ _1321_ _1286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1779__A1 _0852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1520_ _0598_ _0602_ _0603_ _0604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_2_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1451_ net32 _1354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2003_ _1074_ _0976_ _1076_ _1077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_26_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2905_ _0609_ _0567_ _0595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2836_ _0391_ _1407_ _0109_ _0538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1649_ _0672_ _0727_ _0728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1718_ _0795_ _0577_ _0662_ _0796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_53_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2698_ _0052_ _0391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2767_ _1364_ _0323_ _0321_ _0465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_67_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2725__A3 _0259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1503_ _0468_ _0479_ _0489_ _0500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_2483_ _0115_ _0128_ _0151_ _0160_ _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2552_ _0160_ _0151_ _0128_ _0115_ _0236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_2_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2621_ _0244_ _0256_ _0309_ _0310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XTAP_TAPCELL_ROW_38_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2101__A1 _0928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2819_ _0380_ _0519_ _0520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2404__A2 _0073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1921__A4 _0950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2331__A1 _1406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1983_ _1049_ _1052_ _1053_ _1058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2604_ _0284_ _1429_ _0287_ _0290_ _0291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_61_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2466_ _1306_ _1433_ _1287_ _0142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_2535_ _1389_ _0213_ _0216_ _0217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__2322__A1 _1277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2397_ _0064_ _0065_ _1367_ _0066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_6_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2251_ p_shaping_I.counter\[1\] _1323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2320_ _1382_ _1398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_20_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1658__A3 _0693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2182_ _1198_ _1250_ _1251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_18_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1966_ _0909_ _1037_ _1040_ _1041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_28_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1897_ _0967_ _0970_ _0972_ _0791_ _0754_ _0973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_3_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2449_ _1298_ _1379_ _1366_ _1376_ _0123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_11_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2518_ _0051_ _1403_ _0197_ _1387_ _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_54_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1820_ _0887_ _0888_ _0897_ _0758_ _0898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_57_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1751_ _0828_ _0796_ _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1682_ _0759_ _0760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2773__A1 _0328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1923__B _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2303_ _1379_ _1366_ _1300_ _1380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_2234_ _1281_ _1285_ _1293_ _1297_ _1301_ _1303_ _1304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__2525__A1 _0203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2096_ _0731_ _1151_ _1152_ _1154_ _1168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_2165_ _1144_ _1233_ _1234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_0_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1949_ _1023_ _0892_ _0820_ _0914_ _1024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_0_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_8_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1743__B _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1494__A1 _0308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1803_ _0878_ _0880_ _0881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_53_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2921_ _0017_ net56 clknet_1_0__leaf_CLK net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_25_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2783_ _0482_ net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2852_ _0526_ _0545_ _0555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1665_ _0742_ _0743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1596_ net52 _0675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1734_ _0707_ _0812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2746__A1 _0133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1721__A2 _0798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_37_Left_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2217_ _1284_ _1285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_48_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_46_Left_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2079_ _1144_ _1147_ _1152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2148_ _1179_ _1216_ _1217_ _1122_ _1218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_36_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1960__A2 _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_55_Left_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_64_Left_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1450_ _1332_ _1343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2900__A1 _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2002_ _1075_ _0781_ _0602_ _1076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2904_ _0022_ _0594_ _0021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_33_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2835_ _0523_ _0526_ _0537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2766_ _0462_ _0463_ _0464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1648_ _0700_ _0726_ _0727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1579_ _0468_ _0629_ _0599_ _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1717_ _0447_ _0795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2697_ _0380_ _0389_ _0390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_36_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1697__A1 _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2894__B1 _0663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_30_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2620_ _0303_ _0307_ _0309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1502_ _0361_ _0489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_23_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2551_ _0234_ _0165_ _0164_ _0163_ _0235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2482_ _0152_ _0156_ _0159_ _0160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_10_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_38_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2762__B _1390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2818_ _0462_ _1429_ _0501_ _0519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2749_ _0437_ _0445_ _0446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__1679__A1 _0755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2002__B _0602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2391__C _0059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2331__A2 _1301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1982_ _1056_ _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_23_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2601__I _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2603_ _0288_ _0289_ _0290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2534_ _0116_ _0214_ _0215_ _0216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2322__A2 _1399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2396_ _1311_ _0027_ _0065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2465_ _0072_ _0031_ _0106_ _0141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_64_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2561__A2 _1439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1571__B _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2667__B _0025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2250_ _1320_ _1322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_20_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2181_ _1249_ _1221_ _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1500__I _0318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1965_ _0887_ _1039_ _1040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1896_ _0971_ _0855_ _0972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2517_ _0031_ _1368_ _0197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_45_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2448_ _1380_ _0120_ _0121_ _0122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_3_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2379_ _1378_ _0046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_54_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2397__B _1367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1750_ _0733_ _0828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_37_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1681_ _0627_ _0759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_29_Left_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2164_ _1227_ _0734_ _1182_ _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2302_ _1282_ _1379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2233_ _1302_ _1303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_0_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2095_ _1116_ _1119_ _1158_ _1166_ _1167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_51_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2461__A1 _1333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1879_ _0669_ _0924_ _0954_ _0955_ _0956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
X_1948_ _0853_ _1023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_43_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2507__A2 _0073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2920_ _0016_ net56 clknet_1_0__leaf_CLK net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_57_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1733_ _0790_ _0642_ _0810_ _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1802_ _0605_ _0879_ _0880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_31_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2782_ _0477_ _0481_ _0482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2851_ _0554_ net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1595_ _0673_ _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_1664_ _0691_ _0742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_56_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2147_ _1144_ _1216_ _1217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2216_ _1282_ _1283_ _0091_ _1284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_63_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2078_ _1142_ _1143_ _1149_ _1151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_36_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1844__B _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1951__A3 _0636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2001_ _0818_ _1075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2900__A2 _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2903_ _1122_ p_shaping_Q.counter\[0\] _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1716_ _0792_ _0756_ _0793_ _0794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_41_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2834_ _0518_ _0522_ _0536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2765_ _0273_ _0418_ _0463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2696_ _0121_ _0336_ _0388_ _0389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1647_ _0702_ _0725_ _0726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1578_ _0638_ _0654_ _0656_ _0657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_6_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_16_Left_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2407__A1 _0039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2894__A1 _0647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1749__B _0732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2550_ _0166_ _0234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_12_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1501_ _0286_ _0479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_50_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2481_ _0158_ _0159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_58_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_46_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2748_ _0438_ _0444_ _0445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2817_ _0025_ _0517_ _0518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2679_ _0285_ _0370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_1_Left_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1981_ _0617_ _1045_ _1055_ _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_23_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2398__A3 _0037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2533_ _0199_ _0209_ _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2602_ _0168_ _0065_ _0289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_48_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2395_ _1296_ _1313_ _0064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2464_ _0108_ _0140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_57_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1521__A1 _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2234__C1 _1301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2180_ _1168_ _1196_ _1249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1895_ _0665_ _0971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_43_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1964_ _0812_ _0968_ _1038_ _1039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_31_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2447_ _1419_ _0121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2516_ _0194_ _0195_ _0141_ _0101_ _0196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__1898__I _0732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2378_ _0042_ _0044_ _1349_ _0045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_66_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_62_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2790__I0 _0611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_4_Left_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1680_ _0723_ _0758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_29_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2301_ _1346_ _1378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2588__B _1281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2163_ _0022_ _1231_ _1232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2232_ _0157_ _0047_ _1302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2289__A2 _1361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_51_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2094_ _1071_ _1114_ _1166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_0_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2461__A2 _0136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1878_ _0788_ _0941_ _0953_ _0955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1947_ _1020_ _1021_ _1022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_43_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2929__D p_shaping_I.bit_in_1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1660__B1 _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2680__C _0370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_30_Left_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2850_ _0549_ _0552_ _0554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2691__A2 _0033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1663_ _0739_ _0740_ _0659_ _0741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1732_ _0625_ _0810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_40_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1801_ _0619_ _0620_ _0879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2781_ _0407_ _0412_ _0448_ _0478_ _0480_ _0481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_0_13_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1506__I net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1594_ net40 _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_0_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2077_ _1142_ _1143_ _1148_ _0925_ _1149_ _1150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_2146_ _1182_ _1215_ _1216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2215_ _1354_ _1283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_36_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2000_ _1025_ _1074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2902_ _1202_ _0775_ _0587_ _0593_ _0020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2833_ _0535_ net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1715_ _0592_ _0793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1646_ _0705_ _0724_ _0725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1927__A1 _0739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2764_ _0368_ _0462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2695_ _0381_ _0387_ _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1577_ _0655_ _0656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2129_ _0731_ _1178_ _1186_ _1200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_49_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2343__A1 _1422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2915__CLK clknet_1_0__leaf_CLK vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2646__A2 _0203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1500_ _0318_ _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_50_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2480_ _0265_ _0147_ _0158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2885__A2 _1422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2637__A2 _0221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2816_ _0515_ _0516_ _0517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_18_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1629_ _0633_ _0708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2678_ _1359_ _0369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_5_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2747_ _0289_ _0439_ _0443_ _0375_ _0444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2876__A2 _1361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1980_ _0909_ _1048_ _1054_ p_shaping_Q.bit_in_1 _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_23_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2532_ _1345_ _1426_ _0127_ _0214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2601_ _0174_ _0288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_11_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2463_ _0096_ _0138_ _0139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2394_ _0062_ _0063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1818__B1 _0797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout42_I net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwire45 _0299_ net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2794__A1 _0096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1588__A2 _0666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1894_ _0968_ _0969_ _0970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1963_ _0707_ _0763_ _1038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__2528__A1 _0184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2446_ _1298_ _1379_ _1438_ _0031_ _0120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2515_ _1401_ _1312_ _0195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_3_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2377_ _0043_ _0044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_62_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2767__A1 _1364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2519__A1 _0121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2231_ _1298_ _1300_ _1284_ _1301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_0_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2300_ _1374_ _1375_ _1369_ _1377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_2093_ _1162_ _1164_ _1165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2162_ _1229_ _1230_ _1231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_48_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1877_ _0925_ _0941_ _0953_ _0954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1946_ _0672_ _0984_ _1010_ _1011_ _1021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__1972__A2 _0911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2429_ _1331_ _0101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_66_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1963__A2 _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1612__I net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1479__A1 _1397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1800_ _0873_ _0877_ _0878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_57_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1662_ _0626_ _0740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_53_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1731_ _0735_ _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_31_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2780_ _0415_ _0446_ _0480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__1706__A2 _0777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1593_ _0671_ _0672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2214_ net55 _1282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2076_ _1094_ _0998_ _1149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_2145_ _1204_ _1136_ _1078_ _1215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_63_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1642__A1 _0687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1929_ _0806_ _0890_ _1005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1860__C _0719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2370__A2 _1417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1588__B _0553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_33_Left_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_42_Left_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2901_ _1202_ _0590_ _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2832_ _0529_ _0534_ _0535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2763_ _0350_ _0459_ _0460_ _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1576_ _0521_ _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_67_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1645_ _0706_ _0715_ _0718_ _0722_ _0723_ _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_1714_ _0790_ _0778_ _0791_ _0644_ _0792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_41_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2694_ _0383_ _0384_ _0385_ _0386_ _0387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_67_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2128_ _1198_ _1199_ net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2059_ _1125_ _1128_ _1130_ _1131_ _1132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_36_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2343__A2 _1325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2022__A1 _0666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2270__A1 _1330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2746_ _0133_ _0442_ _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2815_ _0148_ _0279_ _0516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1559_ _0631_ _0636_ _0637_ _0638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1628_ _0682_ _0707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2677_ _0288_ _0368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1710__I p_shaping_Q.counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2564__A2 _0033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1620__I _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2600_ _1399_ _0205_ _0037_ _0285_ _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_48_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2393_ p_shaping_I.bit_in_1 _0062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2531_ _0193_ _0210_ _0212_ _0213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2462_ _0072_ _1292_ _1369_ _0138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_64_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwire46 _1100_ net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2729_ _0197_ _0418_ _0424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__2794__A2 _0273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1521__A3 _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2234__A1 _1281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2537__A2 _0044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_56_Right_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1962_ _0807_ _1035_ _1036_ _1037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_50_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1893_ _0943_ _0969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_65_Right_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2445_ _0051_ _0105_ _1341_ _0119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2376_ _1305_ _1336_ _1283_ _0043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2700__A2 _0136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2514_ _1287_ _1290_ _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_54_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2207__B2 _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_2_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2230_ _0058_ _1300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_29_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2092_ _1159_ _1163_ _1164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2161_ _1104_ _1057_ _1230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2694__A1 _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1945_ _0730_ _1009_ _0995_ _0996_ _1020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_28_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1876_ _0951_ _0952_ _0953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_3_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2359_ _1438_ _1439_ _1440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2428_ _1294_ _0100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1660__A2 _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2437__A1 _0105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2676__A1 _0328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1661_ _0329_ _0739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1592_ _0670_ _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1730_ _0807_ _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_40_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2600__A1 _1399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2144_ _1094_ _1213_ _1177_ _0022_ _1214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2213_ _1280_ _1281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2075_ _1144_ _1147_ _1148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1928_ _0735_ _0636_ _1004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1859_ _0810_ _0642_ _0935_ _0936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_31_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_10_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2649__A1 _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1872__A2 _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2900_ _0889_ _0653_ _0589_ _0591_ _0019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1713_ _0297_ _0600_ _0791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_38_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2831_ _0530_ _0533_ _0534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2762_ _0350_ _0432_ _1390_ _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1644_ _0569_ _0723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1575_ _0639_ _0646_ _0650_ _0653_ _0654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2888__B2 _0486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2693_ _0324_ _1416_ _0384_ _0383_ _0385_ _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2127_ _1197_ _1165_ _1167_ _1199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA_fanout65_I net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2058_ _0604_ _1131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_24_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_32_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1854__A2 _0911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1606__A2 _0684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2022__A2 _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2745_ _0440_ _1416_ _0441_ _0442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2814_ _0109_ _0337_ _0514_ _0374_ _0515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2676_ _0328_ _0330_ _0094_ _0367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_14_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1627_ _0542_ _0706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1558_ _0457_ _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1489_ _0340_ _0351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_61_Left_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2261__A2 _1333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2013__A2 _0732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2530_ _1344_ _1425_ _0127_ _0212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_2_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1763__A1 _0752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2392_ _1428_ _0030_ _0041_ _0060_ _0061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_2461_ _1333_ _0136_ _0137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_58_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2798__B _0440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2659_ _0148_ _0350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2728_ _0062_ _0343_ _0342_ _0423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_1_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2234__A2 _1285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_5_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1961_ _0690_ _0989_ _0842_ _1036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_50_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1892_ _0818_ _0653_ _0968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_28_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2513_ _0192_ _0193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2444_ _1314_ _1338_ _1415_ _0101_ _0118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_11_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2375_ _1311_ _1337_ _0042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1672__C2 _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2160_ _1125_ _1227_ _1039_ _1228_ _1229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2091_ _1124_ _1154_ _1155_ _1163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_45_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1944_ _1019_ net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1875_ _0864_ _0878_ _0616_ _0952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_9_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2427_ _0096_ _0032_ _0098_ _0099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_67_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2289_ _1359_ _1361_ _1363_ _1364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2358_ _1353_ _1295_ _1439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_62_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1645__B1 _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2373__A1 _0039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_8_Left_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1660_ _0733_ _0734_ _0736_ _0737_ _0738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_1591_ _0669_ _0670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_33_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2143_ _0671_ _0022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2212_ _1408_ _1280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_63_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2074_ _1078_ _1145_ _1146_ _0771_ _1147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_1858_ _0468_ _0489_ _0691_ _0935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1927_ _0739_ _0703_ _1003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1789_ _0634_ _0382_ _0681_ _0867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_27_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_35_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2897__A2 _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2830_ _0477_ _0481_ _0531_ _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1643_ _0719_ _0721_ _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1712_ _0692_ _0790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_41_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2692_ _0105_ _0221_ _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2761_ _0063_ _0423_ _0458_ _0459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2585__A1 _0234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1574_ _0652_ _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2888__A2 _0133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2126_ _1165_ _1167_ _1197_ _1198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2057_ _1129_ _0969_ _1130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1615__A3 _0693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_24_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2500__A1 _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output39_I net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_38_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2813_ _0285_ _1407_ _0325_ _0514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1626_ _0703_ _0674_ _0704_ _0655_ _0705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_41_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2744_ _0391_ _0203_ _0204_ _0441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2675_ _0347_ _0365_ _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_14_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1557_ _0634_ _0479_ _0635_ _0636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_1488_ net50 _0340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2109_ _1027_ _1180_ _1181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1772__A2 _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2788__A1 _0486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_21_Left_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2460_ _1417_ _1358_ _0136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_48_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2391_ _0045_ _0050_ _0057_ _0059_ _0060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_46_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1609_ _0634_ _0681_ _0688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2589_ _1281_ _0138_ _0273_ _0275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2727_ _0380_ _0421_ _0422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2658_ _0608_ _0342_ _0343_ _0349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_57_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1690__A1 _0754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2473__A3 _0060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1891_ _0743_ _0967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1960_ _0601_ _0736_ _0694_ _1035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1736__A2 _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2443_ _1345_ _1426_ _0116_ _0117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_11_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2512_ _0116_ _0192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2374_ _0035_ _0038_ _1398_ _0040_ _0041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_66_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1672__A1 _0732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1975__A2 _0742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1663__A1 _0739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2090_ _1157_ _1162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_29_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1798__B _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1943_ _1014_ _1018_ _1019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1874_ _0942_ _0945_ _0950_ _0951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_56_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1980__C p_shaping_Q.bit_in_1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_24_Left_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2382__A2 _0048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2426_ _0055_ _0097_ _0098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_67_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1645__A1 _0706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2357_ _1288_ _1438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2288_ _1362_ _1363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_59_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1727__I _0705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1884__A1 _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1590_ p_shaping_Q.counter\[1\] p_shaping_Q.counter\[0\] _0669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_56_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2073_ _0867_ _0849_ _1027_ _1146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2142_ _0618_ _1211_ _1212_ _1213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2211_ _1278_ _1279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_56_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1788_ _0625_ _0759_ _0677_ _0866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1857_ _0795_ _0932_ _0933_ _0851_ _0934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1926_ _0717_ _0679_ _1002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1866__A1 _0687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2409_ _0077_ _0078_ _1371_ _0079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__1618__A1 _0318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2897__A3 _0566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1642_ _0687_ _0704_ _0720_ _0721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1711_ p_shaping_Q.bit_in_2 _0789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_53_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2691_ _0046_ _0033_ _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2760_ _0368_ _1285_ _0073_ _0456_ _0458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_67_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1573_ _0651_ _0640_ _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_6_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2056_ _1079_ _1129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2125_ _1168_ _1196_ _1197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1909_ _0789_ _0985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_32_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2576__A2 _0259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2889_ _0486_ _0581_ _0584_ _0014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_4_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1839__A1 _0818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput4 net4 I[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__2520__B _0101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2007__A1 _0887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2812_ _0513_ net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2743_ _1372_ _0440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1625_ _0676_ _0704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1556_ _0414_ _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2674_ _0332_ _0354_ _0365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1487_ _0318_ _0329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2039_ _1107_ _1111_ _1082_ _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2108_ _0689_ _1023_ _1180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1735__I _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2788__A2 _0080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2390_ _1316_ _0059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2726_ _0368_ _0419_ _0420_ _0283_ _0421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_6_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1608_ _0600_ _0687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1539_ _0612_ _0619_ _0620_ _0621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2703__A2 _1340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2588_ _0138_ _0273_ _1281_ _0274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2657_ _0333_ _0341_ _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_40_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_5_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1890_ _0965_ _0956_ _0966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1736__A3 _0755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2442_ p_shaping_I.bit_in_2 _0116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2373_ _0039_ _0113_ _1317_ _0040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2511_ _0187_ _0190_ _0191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_49_Left_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1975__A3 _0693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2709_ _0115_ _0390_ _0401_ _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_58_Left_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_2_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_67_Left_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_61_Right_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1718__A3 _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1942_ _1015_ _1017_ _1018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1873_ _0946_ _0947_ _0949_ _0770_ _0950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_43_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1590__A1 p_shaping_Q.counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2356_ _1401_ _1303_ _1308_ _1437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__2382__A3 _0049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2425_ _1356_ _1303_ _0097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_67_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2287_ _1288_ _1362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_62_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1636__A2 _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1918__I _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2210_ _0135_ _1278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_56_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2072_ _1086_ _0847_ _1137_ _1145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_2141_ _1109_ _1211_ _1212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_56_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1925_ _0807_ _0734_ _0999_ _1000_ _1001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_44_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1787_ _0863_ _0864_ _0865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1856_ _0790_ _0810_ _0778_ _0933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_31_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2339_ _1292_ _1415_ _1416_ _1417_ _1418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_2408_ _1402_ _1307_ _1362_ _0078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_27_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2034__A2 _1092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1641_ _0447_ _0720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_1710_ p_shaping_Q.counter\[1\] _0788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1793__A1 _0308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1572_ _0632_ _0651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_21_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2690_ _0182_ _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2124_ _1188_ _1195_ _1196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2055_ _1126_ _1127_ _1087_ _0874_ _1128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__1558__I _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1839_ _0818_ _0704_ _0916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1908_ _0980_ _0983_ _0984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_44_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2888_ _0583_ _0133_ _0581_ _0486_ _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_4_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1468__I net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput5 net5 I[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput40 net40 addQ[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__2327__I0 _1314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2299__I _1337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_1_0__f_CLK clknet_0_CLK clknet_1_0__leaf_CLK vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__2255__A2 _1325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2007__A2 _1049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2811_ _0485_ _0508_ _0512_ _0513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2742_ _0375_ _1422_ _0439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1624_ _0664_ _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1555_ _0633_ _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2673_ _0364_ net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2107_ _0804_ _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1486_ net51 _0318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_fanout63_I net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2038_ _1082_ _1107_ _1111_ _1112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_49_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2228__A2 _1296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2725_ _0284_ _0294_ _0259_ _0420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_6_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2656_ _0333_ _0341_ _0345_ _0305_ _0346_ _0347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_1607_ _0521_ _0680_ _0683_ _0685_ _0686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__1911__A1 _0694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1538_ net62 p_shaping_Q.ctl_1 _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1469_ net35 _0135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2587_ _1310_ _1338_ _0273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__1520__B _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1978__A1 _0719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1656__I _0684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2510_ _0188_ _0111_ _0610_ _0190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2372_ _1326_ _0039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_11_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2441_ _1324_ _0115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_59_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2639_ _0283_ _0322_ _0327_ _0328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_6_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2708_ _0115_ _0390_ _0401_ _0402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_65_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1941_ _0837_ _0904_ _1016_ _0962_ _1017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_56_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1872_ _0795_ _0811_ _0948_ _0949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_16_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2424_ _1278_ _1280_ _0096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_2355_ _1306_ _1287_ _1290_ _1436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2286_ _1360_ _1361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_59_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_13_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2140_ _1125_ _1192_ _1210_ _1211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2521__A1 _0039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2071_ _1083_ _1144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_29_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1855_ _0869_ _0687_ _0932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1924_ _0761_ _0943_ _0842_ _1000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_8_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1786_ _0758_ _0776_ _0784_ _0700_ _0864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_31_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2269_ _1337_ _1339_ _1340_ _1308_ _1341_ _1342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_2338_ _1336_ _1417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2407_ _0039_ _0076_ _0077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_67_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1857__A3 _0933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1640_ _0532_ _0719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1571_ _0647_ _0649_ _0645_ _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__1793__A2 _0720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2123_ _1194_ _1195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_49_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2054_ _1038_ _0968_ _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1838_ _0914_ _0813_ _0915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1907_ _0752_ _0982_ _0983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2887_ _0582_ _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1769_ _0649_ _0652_ _0847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_40_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput41 net41 addQ[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__1775__A2 _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput30 net55 addI[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_23_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput6 net6 I[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_46_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2810_ _0509_ _0510_ _0512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2741_ _0367_ _0438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2672_ _0356_ _0363_ _0364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1623_ _0701_ _0702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1485_ _0297_ _0308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1554_ _0632_ _0633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_1_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
.ends

